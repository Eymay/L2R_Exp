`timescale 1ns / 1ps
module L2RExp (Done,
    clk,
    rst,
    start,
    A,
    B,
    C);
 output Done;
 input clk;
 input rst;
 input start;
 input [15:0] A;
 input [15:0] B;
 output [31:0] C;

 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire clknet_0_clk;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire \control_unit.LoadA ;
 wire \control_unit.LoadC ;
 wire \control_unit.LoadCoun ;
 wire \control_unit.S_C[0] ;
 wire \control_unit.S_C[1] ;
 wire \control_unit.S_Coun ;
 wire \control_unit.ShiftB ;
 wire \control_unit.regBk ;
 wire \control_unit.state[0] ;
 wire \control_unit.state[1] ;
 wire \control_unit.state[2] ;
 wire \datapath.Counter[0] ;
 wire \datapath.Counter[1] ;
 wire \datapath.Counter[2] ;
 wire \datapath.Counter[3] ;
 wire \datapath.Counter[4] ;
 wire \datapath.MultiplierAC.PPG0.X[0] ;
 wire \datapath.MultiplierAC.PPG0.X[10] ;
 wire \datapath.MultiplierAC.PPG0.X[11] ;
 wire \datapath.MultiplierAC.PPG0.X[12] ;
 wire \datapath.MultiplierAC.PPG0.X[13] ;
 wire \datapath.MultiplierAC.PPG0.X[14] ;
 wire \datapath.MultiplierAC.PPG0.X[15] ;
 wire \datapath.MultiplierAC.PPG0.X[1] ;
 wire \datapath.MultiplierAC.PPG0.X[2] ;
 wire \datapath.MultiplierAC.PPG0.X[3] ;
 wire \datapath.MultiplierAC.PPG0.X[4] ;
 wire \datapath.MultiplierAC.PPG0.X[5] ;
 wire \datapath.MultiplierAC.PPG0.X[6] ;
 wire \datapath.MultiplierAC.PPG0.X[7] ;
 wire \datapath.MultiplierAC.PPG0.X[8] ;
 wire \datapath.MultiplierAC.PPG0.X[9] ;
 wire \datapath.MultiplierAC.PPG0.Y[0] ;
 wire \datapath.MultiplierAC.PPG0.Y[10] ;
 wire \datapath.MultiplierAC.PPG0.Y[11] ;
 wire \datapath.MultiplierAC.PPG0.Y[12] ;
 wire \datapath.MultiplierAC.PPG0.Y[13] ;
 wire \datapath.MultiplierAC.PPG0.Y[14] ;
 wire \datapath.MultiplierAC.PPG0.Y[15] ;
 wire \datapath.MultiplierAC.PPG0.Y[1] ;
 wire \datapath.MultiplierAC.PPG0.Y[2] ;
 wire \datapath.MultiplierAC.PPG0.Y[3] ;
 wire \datapath.MultiplierAC.PPG0.Y[4] ;
 wire \datapath.MultiplierAC.PPG0.Y[5] ;
 wire \datapath.MultiplierAC.PPG0.Y[6] ;
 wire \datapath.MultiplierAC.PPG0.Y[7] ;
 wire \datapath.MultiplierAC.PPG0.Y[8] ;
 wire \datapath.MultiplierAC.PPG0.Y[9] ;
 wire \datapath.RegB[0] ;
 wire \datapath.RegB[10] ;
 wire \datapath.RegB[11] ;
 wire \datapath.RegB[12] ;
 wire \datapath.RegB[13] ;
 wire \datapath.RegB[14] ;
 wire \datapath.RegB[1] ;
 wire \datapath.RegB[2] ;
 wire \datapath.RegB[3] ;
 wire \datapath.RegB[4] ;
 wire \datapath.RegB[5] ;
 wire \datapath.RegB[6] ;
 wire \datapath.RegB[7] ;
 wire \datapath.RegB[8] ;
 wire \datapath.RegB[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0__1442_;
 wire clknet_1_0__leaf__1442_;
 wire clknet_1_1__leaf__1442_;

 sky130_fd_sc_hd__inv_2 _2194_ (.A(\control_unit.LoadA ),
    .Y(_1045_));
 sky130_fd_sc_hd__buf_4 _2195_ (.A(_1045_),
    .X(_1056_));
 sky130_fd_sc_hd__clkbuf_4 _2196_ (.A(net33),
    .X(_1067_));
 sky130_fd_sc_hd__buf_4 _2197_ (.A(_1067_),
    .X(_1078_));
 sky130_fd_sc_hd__clkbuf_8 _2198_ (.A(\control_unit.LoadA ),
    .X(_1089_));
 sky130_fd_sc_hd__or2_1 _2199_ (.A(\datapath.MultiplierAC.PPG0.Y[15] ),
    .B(_1089_),
    .X(_1100_));
 sky130_fd_sc_hd__o211a_1 _2200_ (.A1(net7),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1100_),
    .X(_0074_));
 sky130_fd_sc_hd__inv_2 _2201_ (.A(\datapath.MultiplierAC.PPG0.Y[14] ),
    .Y(_1121_));
 sky130_fd_sc_hd__nand2_1 _2202_ (.A(_1056_),
    .B(_1121_),
    .Y(_1132_));
 sky130_fd_sc_hd__o211a_1 _2203_ (.A1(net6),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1132_),
    .X(_0073_));
 sky130_fd_sc_hd__or2_1 _2204_ (.A(_1089_),
    .B(\datapath.MultiplierAC.PPG0.Y[13] ),
    .X(_1153_));
 sky130_fd_sc_hd__o211a_1 _2205_ (.A1(net5),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1153_),
    .X(_0072_));
 sky130_fd_sc_hd__or2_1 _2206_ (.A(_1089_),
    .B(\datapath.MultiplierAC.PPG0.Y[12] ),
    .X(_1173_));
 sky130_fd_sc_hd__o211a_1 _2207_ (.A1(net4),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1173_),
    .X(_0071_));
 sky130_fd_sc_hd__inv_2 _2208_ (.A(\datapath.MultiplierAC.PPG0.Y[11] ),
    .Y(_1194_));
 sky130_fd_sc_hd__nand2_1 _2209_ (.A(_1056_),
    .B(_1194_),
    .Y(_1205_));
 sky130_fd_sc_hd__o211a_1 _2210_ (.A1(net3),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1205_),
    .X(_0070_));
 sky130_fd_sc_hd__clkbuf_8 _2211_ (.A(_1045_),
    .X(_1226_));
 sky130_fd_sc_hd__inv_2 _2212_ (.A(\datapath.MultiplierAC.PPG0.Y[10] ),
    .Y(_1237_));
 sky130_fd_sc_hd__nand2_1 _2213_ (.A(_1226_),
    .B(_1237_),
    .Y(_1248_));
 sky130_fd_sc_hd__o211a_1 _2214_ (.A1(net2),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1248_),
    .X(_0069_));
 sky130_fd_sc_hd__or2_1 _2215_ (.A(_1089_),
    .B(\datapath.MultiplierAC.PPG0.Y[9] ),
    .X(_1269_));
 sky130_fd_sc_hd__o211a_1 _2216_ (.A1(net16),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1269_),
    .X(_0068_));
 sky130_fd_sc_hd__or2_1 _2217_ (.A(_1089_),
    .B(\datapath.MultiplierAC.PPG0.Y[8] ),
    .X(_1290_));
 sky130_fd_sc_hd__o211a_1 _2218_ (.A1(net15),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1290_),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_4 _2219_ (.A(\datapath.MultiplierAC.PPG0.Y[7] ),
    .X(_1311_));
 sky130_fd_sc_hd__or2_1 _2220_ (.A(_1089_),
    .B(_1311_),
    .X(_1322_));
 sky130_fd_sc_hd__o211a_1 _2221_ (.A1(net14),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1322_),
    .X(_0066_));
 sky130_fd_sc_hd__clkbuf_4 _2222_ (.A(\datapath.MultiplierAC.PPG0.Y[6] ),
    .X(_1343_));
 sky130_fd_sc_hd__inv_2 _2223_ (.A(_1343_),
    .Y(_1354_));
 sky130_fd_sc_hd__nand2_1 _2224_ (.A(_1226_),
    .B(_1354_),
    .Y(_1364_));
 sky130_fd_sc_hd__o211a_1 _2225_ (.A1(net13),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1364_),
    .X(_0065_));
 sky130_fd_sc_hd__buf_4 _2226_ (.A(\datapath.MultiplierAC.PPG0.Y[5] ),
    .X(_1379_));
 sky130_fd_sc_hd__inv_2 _2227_ (.A(_1379_),
    .Y(_1387_));
 sky130_fd_sc_hd__nand2_1 _2228_ (.A(_1226_),
    .B(_1387_),
    .Y(_1395_));
 sky130_fd_sc_hd__o211a_1 _2229_ (.A1(net12),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1395_),
    .X(_0064_));
 sky130_fd_sc_hd__buf_4 _2230_ (.A(\datapath.MultiplierAC.PPG0.Y[4] ),
    .X(_1411_));
 sky130_fd_sc_hd__or2_1 _2231_ (.A(_1089_),
    .B(_1411_),
    .X(_1419_));
 sky130_fd_sc_hd__o211a_1 _2232_ (.A1(net11),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1419_),
    .X(_0063_));
 sky130_fd_sc_hd__buf_4 _2233_ (.A(\datapath.MultiplierAC.PPG0.Y[3] ),
    .X(_1435_));
 sky130_fd_sc_hd__or2_1 _2234_ (.A(_1089_),
    .B(_1435_),
    .X(_1443_));
 sky130_fd_sc_hd__o211a_1 _2235_ (.A1(net10),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1443_),
    .X(_0062_));
 sky130_fd_sc_hd__buf_4 _2236_ (.A(\datapath.MultiplierAC.PPG0.Y[2] ),
    .X(_1448_));
 sky130_fd_sc_hd__inv_2 _2237_ (.A(_1448_),
    .Y(_1457_));
 sky130_fd_sc_hd__nand2_1 _2238_ (.A(_1226_),
    .B(_1457_),
    .Y(_1462_));
 sky130_fd_sc_hd__o211a_1 _2239_ (.A1(net9),
    .A2(_1056_),
    .B1(_1078_),
    .C1(_1462_),
    .X(_0061_));
 sky130_fd_sc_hd__buf_8 _2240_ (.A(\datapath.MultiplierAC.PPG0.Y[1] ),
    .X(_1463_));
 sky130_fd_sc_hd__inv_2 _2241_ (.A(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__nand2_1 _2242_ (.A(_1226_),
    .B(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__o211a_1 _2243_ (.A1(net8),
    .A2(_1056_),
    .B1(_1067_),
    .C1(_1465_),
    .X(_0060_));
 sky130_fd_sc_hd__buf_8 _2244_ (.A(\datapath.MultiplierAC.PPG0.Y[0] ),
    .X(_1466_));
 sky130_fd_sc_hd__or2_1 _2245_ (.A(_1089_),
    .B(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__o211a_1 _2246_ (.A1(net1),
    .A2(_1056_),
    .B1(_1067_),
    .C1(_1467_),
    .X(_0059_));
 sky130_fd_sc_hd__or4_1 _2247_ (.A(net3),
    .B(net2),
    .C(net16),
    .D(net15),
    .X(_1468_));
 sky130_fd_sc_hd__or4_1 _2248_ (.A(net7),
    .B(net6),
    .C(net5),
    .D(net4),
    .X(_1469_));
 sky130_fd_sc_hd__or4_1 _2249_ (.A(net10),
    .B(net9),
    .C(net8),
    .D(net1),
    .X(_1470_));
 sky130_fd_sc_hd__or4_1 _2250_ (.A(net14),
    .B(net13),
    .C(net12),
    .D(net11),
    .X(_1471_));
 sky130_fd_sc_hd__or4_1 _2251_ (.A(_1468_),
    .B(_1469_),
    .C(_1470_),
    .D(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__buf_6 _2252_ (.A(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__buf_12 _2253_ (.A(\datapath.MultiplierAC.PPG0.X[0] ),
    .X(_1474_));
 sky130_fd_sc_hd__buf_12 _2254_ (.A(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__nor3_1 _2255_ (.A(\datapath.Counter[4] ),
    .B(\datapath.Counter[3] ),
    .C(\datapath.Counter[0] ),
    .Y(_1476_));
 sky130_fd_sc_hd__nor2_1 _2256_ (.A(\datapath.Counter[2] ),
    .B(\datapath.Counter[1] ),
    .Y(_1477_));
 sky130_fd_sc_hd__nand2_2 _2257_ (.A(_1476_),
    .B(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__inv_6 _2258_ (.A(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__and3_1 _2259_ (.A(_1473_),
    .B(_1475_),
    .C(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__clkbuf_1 _2260_ (.A(_1480_),
    .X(net35));
 sky130_fd_sc_hd__buf_12 _2261_ (.A(\datapath.MultiplierAC.PPG0.X[1] ),
    .X(_1481_));
 sky130_fd_sc_hd__buf_8 _2262_ (.A(_1481_),
    .X(_1482_));
 sky130_fd_sc_hd__and3_1 _2263_ (.A(_1473_),
    .B(_1482_),
    .C(_1479_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_1 _2264_ (.A(_1483_),
    .X(net42));
 sky130_fd_sc_hd__buf_8 _2265_ (.A(\datapath.MultiplierAC.PPG0.X[2] ),
    .X(_1484_));
 sky130_fd_sc_hd__buf_8 _2266_ (.A(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__and3_1 _2267_ (.A(_1473_),
    .B(_1485_),
    .C(_1479_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _2268_ (.A(_1486_),
    .X(net43));
 sky130_fd_sc_hd__buf_8 _2269_ (.A(\datapath.MultiplierAC.PPG0.X[3] ),
    .X(_1487_));
 sky130_fd_sc_hd__buf_8 _2270_ (.A(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__and3_1 _2271_ (.A(_1473_),
    .B(_1488_),
    .C(_1479_),
    .X(_1489_));
 sky130_fd_sc_hd__clkbuf_1 _2272_ (.A(_1489_),
    .X(net44));
 sky130_fd_sc_hd__buf_12 _2273_ (.A(\datapath.MultiplierAC.PPG0.X[4] ),
    .X(_1490_));
 sky130_fd_sc_hd__and3_1 _2274_ (.A(_1473_),
    .B(_1490_),
    .C(_1479_),
    .X(_1491_));
 sky130_fd_sc_hd__clkbuf_1 _2275_ (.A(_1491_),
    .X(net45));
 sky130_fd_sc_hd__buf_8 _2276_ (.A(\datapath.MultiplierAC.PPG0.X[5] ),
    .X(_1492_));
 sky130_fd_sc_hd__and3_1 _2277_ (.A(_1473_),
    .B(_1492_),
    .C(_1479_),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_1 _2278_ (.A(_1493_),
    .X(net46));
 sky130_fd_sc_hd__buf_12 _2279_ (.A(\datapath.MultiplierAC.PPG0.X[6] ),
    .X(_1494_));
 sky130_fd_sc_hd__and3_1 _2280_ (.A(_1473_),
    .B(_1494_),
    .C(_1479_),
    .X(_1495_));
 sky130_fd_sc_hd__clkbuf_1 _2281_ (.A(_1495_),
    .X(net47));
 sky130_fd_sc_hd__buf_8 _2282_ (.A(\datapath.MultiplierAC.PPG0.X[7] ),
    .X(_1496_));
 sky130_fd_sc_hd__and3_1 _2283_ (.A(_1473_),
    .B(_1496_),
    .C(_1479_),
    .X(_1497_));
 sky130_fd_sc_hd__clkbuf_1 _2284_ (.A(_1497_),
    .X(net48));
 sky130_fd_sc_hd__buf_6 _2285_ (.A(\datapath.MultiplierAC.PPG0.X[8] ),
    .X(_1498_));
 sky130_fd_sc_hd__and3_1 _2286_ (.A(_1473_),
    .B(_1498_),
    .C(_1479_),
    .X(_1499_));
 sky130_fd_sc_hd__clkbuf_1 _2287_ (.A(_1499_),
    .X(net49));
 sky130_fd_sc_hd__buf_6 _2288_ (.A(\datapath.MultiplierAC.PPG0.X[9] ),
    .X(_1500_));
 sky130_fd_sc_hd__and3_1 _2289_ (.A(_1473_),
    .B(_1500_),
    .C(_1479_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _2290_ (.A(_1501_),
    .X(net50));
 sky130_fd_sc_hd__buf_6 _2291_ (.A(\datapath.MultiplierAC.PPG0.X[10] ),
    .X(_1502_));
 sky130_fd_sc_hd__and3_1 _2292_ (.A(_1473_),
    .B(_1502_),
    .C(_1479_),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_1 _2293_ (.A(_1503_),
    .X(net36));
 sky130_fd_sc_hd__buf_4 _2294_ (.A(\datapath.MultiplierAC.PPG0.X[11] ),
    .X(_1504_));
 sky130_fd_sc_hd__and3_1 _2295_ (.A(_1473_),
    .B(_1504_),
    .C(_1479_),
    .X(_1505_));
 sky130_fd_sc_hd__clkbuf_1 _2296_ (.A(_1505_),
    .X(net37));
 sky130_fd_sc_hd__and3_1 _2297_ (.A(_1473_),
    .B(\datapath.MultiplierAC.PPG0.X[12] ),
    .C(_1479_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_1 _2298_ (.A(_1506_),
    .X(net38));
 sky130_fd_sc_hd__and3_1 _2299_ (.A(_1473_),
    .B(\datapath.MultiplierAC.PPG0.X[13] ),
    .C(_1479_),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_1 _2300_ (.A(_1507_),
    .X(net39));
 sky130_fd_sc_hd__and3_1 _2301_ (.A(_1473_),
    .B(\datapath.MultiplierAC.PPG0.X[14] ),
    .C(_1479_),
    .X(_1508_));
 sky130_fd_sc_hd__clkbuf_1 _2302_ (.A(_1508_),
    .X(net40));
 sky130_fd_sc_hd__and3_1 _2303_ (.A(_1473_),
    .B(\datapath.MultiplierAC.PPG0.X[15] ),
    .C(_1479_),
    .X(_1509_));
 sky130_fd_sc_hd__clkbuf_1 _2304_ (.A(_1509_),
    .X(net41));
 sky130_fd_sc_hd__clkinv_4 _2305_ (.A(_1475_),
    .Y(_1510_));
 sky130_fd_sc_hd__nand2_1 _2306_ (.A(_1510_),
    .B(\control_unit.S_C[0] ),
    .Y(_1511_));
 sky130_fd_sc_hd__clkinv_2 _2307_ (.A(\control_unit.S_C[1] ),
    .Y(_1512_));
 sky130_fd_sc_hd__nor2_8 _2308_ (.A(\control_unit.S_C[0] ),
    .B(_1512_),
    .Y(_1513_));
 sky130_fd_sc_hd__nand2_1 _2309_ (.A(_1466_),
    .B(_1474_),
    .Y(_1514_));
 sky130_fd_sc_hd__inv_2 _2310_ (.A(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__a22o_1 _2311_ (.A1(_1511_),
    .A2(_1512_),
    .B1(_1513_),
    .B2(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__buf_4 _2312_ (.A(\control_unit.LoadC ),
    .X(_1517_));
 sky130_fd_sc_hd__clkinv_4 _2313_ (.A(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hd__a21oi_1 _2314_ (.A1(\control_unit.S_C[0] ),
    .A2(\control_unit.S_C[1] ),
    .B1(_1518_),
    .Y(_1519_));
 sky130_fd_sc_hd__and3_1 _2315_ (.A(_1516_),
    .B(_1067_),
    .C(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_1 _2316_ (.A(_1520_),
    .X(_0016_));
 sky130_fd_sc_hd__nor2_1 _2317_ (.A(_1517_),
    .B(_1510_),
    .Y(_1521_));
 sky130_fd_sc_hd__a22o_1 _2318_ (.A1(_1463_),
    .A2(_1475_),
    .B1(_1466_),
    .B2(_1482_),
    .X(_1522_));
 sky130_fd_sc_hd__nand2_1 _2319_ (.A(_1463_),
    .B(_1481_),
    .Y(_1523_));
 sky130_fd_sc_hd__inv_2 _2320_ (.A(_1523_),
    .Y(_1524_));
 sky130_fd_sc_hd__nand2_1 _2321_ (.A(_1515_),
    .B(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__and4_1 _2322_ (.A(_1522_),
    .B(_1513_),
    .C(_1519_),
    .D(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__o21a_1 _2323_ (.A1(_1521_),
    .A2(_1526_),
    .B1(_1078_),
    .X(_0017_));
 sky130_fd_sc_hd__nand2_2 _2324_ (.A(_1466_),
    .B(_1484_),
    .Y(_1527_));
 sky130_fd_sc_hd__nand2_1 _2325_ (.A(_1524_),
    .B(_1527_),
    .Y(_1528_));
 sky130_fd_sc_hd__inv_2 _2326_ (.A(_1527_),
    .Y(_1529_));
 sky130_fd_sc_hd__nand2_1 _2327_ (.A(_1529_),
    .B(_1523_),
    .Y(_1530_));
 sky130_fd_sc_hd__nand3_1 _2328_ (.A(_1525_),
    .B(_1528_),
    .C(_1530_),
    .Y(_1531_));
 sky130_fd_sc_hd__nand3_1 _2329_ (.A(_1515_),
    .B(_1524_),
    .C(_1527_),
    .Y(_1532_));
 sky130_fd_sc_hd__nand2_1 _2330_ (.A(_1448_),
    .B(_1475_),
    .Y(_1533_));
 sky130_fd_sc_hd__inv_2 _2331_ (.A(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__a21o_1 _2332_ (.A1(_1531_),
    .A2(_1532_),
    .B1(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__nand3_1 _2333_ (.A(_1531_),
    .B(_1534_),
    .C(_1532_),
    .Y(_1536_));
 sky130_fd_sc_hd__clkinv_2 _2334_ (.A(\control_unit.S_C[0] ),
    .Y(_1537_));
 sky130_fd_sc_hd__nor2_8 _2335_ (.A(\control_unit.S_C[1] ),
    .B(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hd__inv_2 _2336_ (.A(_1482_),
    .Y(_1539_));
 sky130_fd_sc_hd__nor2_1 _2337_ (.A(_1475_),
    .B(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__a32o_1 _2338_ (.A1(_1535_),
    .A2(_1513_),
    .A3(_1536_),
    .B1(_1538_),
    .B2(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__nand2_1 _2339_ (.A(_1541_),
    .B(_1517_),
    .Y(_1542_));
 sky130_fd_sc_hd__nand2_1 _2340_ (.A(_1518_),
    .B(_1482_),
    .Y(_1543_));
 sky130_fd_sc_hd__inv_2 _2341_ (.A(_1067_),
    .Y(_1544_));
 sky130_fd_sc_hd__clkbuf_8 _2342_ (.A(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__a21oi_1 _2343_ (.A1(_1542_),
    .A2(_1543_),
    .B1(_1545_),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2_1 _2344_ (.A(_1435_),
    .B(_1475_),
    .Y(_1546_));
 sky130_fd_sc_hd__a21oi_1 _2345_ (.A1(_1514_),
    .A2(_1527_),
    .B1(_1523_),
    .Y(_1547_));
 sky130_fd_sc_hd__inv_2 _2346_ (.A(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__nand2_1 _2347_ (.A(_1463_),
    .B(_1487_),
    .Y(_1549_));
 sky130_fd_sc_hd__nor2_1 _2348_ (.A(_1527_),
    .B(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__inv_2 _2349_ (.A(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__nand2_1 _2350_ (.A(_1463_),
    .B(_1484_),
    .Y(_1552_));
 sky130_fd_sc_hd__nand2_1 _2351_ (.A(_1466_),
    .B(_1487_),
    .Y(_1553_));
 sky130_fd_sc_hd__nand2_1 _2352_ (.A(_1552_),
    .B(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__nand2_1 _2353_ (.A(_1551_),
    .B(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__nand2_1 _2354_ (.A(_1548_),
    .B(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__inv_2 _2355_ (.A(_1554_),
    .Y(_1557_));
 sky130_fd_sc_hd__nor2_1 _2356_ (.A(_1550_),
    .B(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__nand2_1 _2357_ (.A(_1558_),
    .B(_1547_),
    .Y(_1559_));
 sky130_fd_sc_hd__nand2_1 _2358_ (.A(_1556_),
    .B(_1559_),
    .Y(_1560_));
 sky130_fd_sc_hd__nand2_1 _2359_ (.A(_1448_),
    .B(_1482_),
    .Y(_1561_));
 sky130_fd_sc_hd__nand2_1 _2360_ (.A(_1560_),
    .B(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__nand3b_1 _2361_ (.A_N(_1561_),
    .B(_1556_),
    .C(_1559_),
    .Y(_1563_));
 sky130_fd_sc_hd__inv_2 _2362_ (.A(_1536_),
    .Y(_1564_));
 sky130_fd_sc_hd__a21o_1 _2363_ (.A1(_1562_),
    .A2(_1563_),
    .B1(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__nand3_1 _2364_ (.A(_1562_),
    .B(_1563_),
    .C(_1564_),
    .Y(_1566_));
 sky130_fd_sc_hd__nand2_1 _2365_ (.A(_1565_),
    .B(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__nor2_1 _2366_ (.A(_1546_),
    .B(_1567_),
    .Y(_1568_));
 sky130_fd_sc_hd__inv_2 _2367_ (.A(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__nand2_1 _2368_ (.A(_1567_),
    .B(_1546_),
    .Y(_1570_));
 sky130_fd_sc_hd__nand2_1 _2369_ (.A(_1488_),
    .B(_1475_),
    .Y(_1571_));
 sky130_fd_sc_hd__nand2_2 _2370_ (.A(_1484_),
    .B(_1481_),
    .Y(_1572_));
 sky130_fd_sc_hd__nand2_1 _2371_ (.A(_1571_),
    .B(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__nand2_4 _2372_ (.A(_1481_),
    .B(_1474_),
    .Y(_1574_));
 sky130_fd_sc_hd__clkinv_4 _2373_ (.A(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hd__nand2_2 _2374_ (.A(_1487_),
    .B(_1484_),
    .Y(_1576_));
 sky130_fd_sc_hd__nand3_1 _2375_ (.A(_1573_),
    .B(_1575_),
    .C(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__nand3_1 _2376_ (.A(_1571_),
    .B(_1572_),
    .C(_1574_),
    .Y(_1578_));
 sky130_fd_sc_hd__nand2_1 _2377_ (.A(_1577_),
    .B(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__nand2_1 _2378_ (.A(_1579_),
    .B(_1572_),
    .Y(_1580_));
 sky130_fd_sc_hd__inv_2 _2379_ (.A(_1571_),
    .Y(_1581_));
 sky130_fd_sc_hd__inv_2 _2380_ (.A(_1572_),
    .Y(_1582_));
 sky130_fd_sc_hd__o21ai_1 _2381_ (.A1(_1574_),
    .A2(_1581_),
    .B1(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__nand2_1 _2382_ (.A(_1485_),
    .B(_1475_),
    .Y(_1584_));
 sky130_fd_sc_hd__inv_2 _2383_ (.A(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__a21o_1 _2384_ (.A1(_1580_),
    .A2(_1583_),
    .B1(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__o2111ai_2 _2385_ (.A1(_1539_),
    .A2(_1576_),
    .B1(_1485_),
    .C1(_1475_),
    .D1(_1573_),
    .Y(_1587_));
 sky130_fd_sc_hd__a21o_1 _2386_ (.A1(_1586_),
    .A2(_1587_),
    .B1(_1581_),
    .X(_1588_));
 sky130_fd_sc_hd__nand3_1 _2387_ (.A(_1586_),
    .B(_1581_),
    .C(_1587_),
    .Y(_1589_));
 sky130_fd_sc_hd__and3_1 _2388_ (.A(_1588_),
    .B(_1589_),
    .C(_1538_),
    .X(_1590_));
 sky130_fd_sc_hd__a31o_1 _2389_ (.A1(_1513_),
    .A2(_1569_),
    .A3(_1570_),
    .B1(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__nand2_1 _2390_ (.A(_1591_),
    .B(_1517_),
    .Y(_1592_));
 sky130_fd_sc_hd__nand2_1 _2391_ (.A(_1518_),
    .B(_1485_),
    .Y(_1593_));
 sky130_fd_sc_hd__a21oi_1 _2392_ (.A1(_1592_),
    .A2(_1593_),
    .B1(_1545_),
    .Y(_0019_));
 sky130_fd_sc_hd__nand2_2 _2393_ (.A(_1411_),
    .B(_1474_),
    .Y(_1594_));
 sky130_fd_sc_hd__nand2_1 _2394_ (.A(_1559_),
    .B(_1551_),
    .Y(_1595_));
 sky130_fd_sc_hd__nand2_1 _2395_ (.A(_1463_),
    .B(_1490_),
    .Y(_1596_));
 sky130_fd_sc_hd__nand2_1 _2396_ (.A(_1466_),
    .B(\datapath.MultiplierAC.PPG0.X[4] ),
    .Y(_1597_));
 sky130_fd_sc_hd__nand2_1 _2397_ (.A(_1549_),
    .B(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__o21ai_1 _2398_ (.A1(_1553_),
    .A2(_1596_),
    .B1(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__inv_2 _2399_ (.A(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__nand2_1 _2400_ (.A(_1595_),
    .B(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__nand2_1 _2401_ (.A(_1448_),
    .B(_1485_),
    .Y(_1602_));
 sky130_fd_sc_hd__inv_2 _2402_ (.A(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__nand3_1 _2403_ (.A(_1559_),
    .B(_1551_),
    .C(_1599_),
    .Y(_1604_));
 sky130_fd_sc_hd__nand3_2 _2404_ (.A(_1601_),
    .B(_1603_),
    .C(_1604_),
    .Y(_1605_));
 sky130_fd_sc_hd__nand2_1 _2405_ (.A(_1595_),
    .B(_1599_),
    .Y(_1606_));
 sky130_fd_sc_hd__nand3_1 _2406_ (.A(_1559_),
    .B(_1551_),
    .C(_1600_),
    .Y(_1607_));
 sky130_fd_sc_hd__nand3_1 _2407_ (.A(_1606_),
    .B(_1602_),
    .C(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__nand2_1 _2408_ (.A(_1605_),
    .B(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__nand3_1 _2409_ (.A(_1609_),
    .B(_1563_),
    .C(_1566_),
    .Y(_1610_));
 sky130_fd_sc_hd__inv_2 _2410_ (.A(_1609_),
    .Y(_1611_));
 sky130_fd_sc_hd__nand2_1 _2411_ (.A(_1566_),
    .B(_1563_),
    .Y(_1612_));
 sky130_fd_sc_hd__nand2_1 _2412_ (.A(_1611_),
    .B(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__nand2_1 _2413_ (.A(_1610_),
    .B(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__nand2_1 _2414_ (.A(_1435_),
    .B(_1482_),
    .Y(_1615_));
 sky130_fd_sc_hd__nand2_1 _2415_ (.A(_1614_),
    .B(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__nand3b_1 _2416_ (.A_N(_1615_),
    .B(_1610_),
    .C(_1613_),
    .Y(_1617_));
 sky130_fd_sc_hd__a21o_1 _2417_ (.A1(_1616_),
    .A2(_1617_),
    .B1(_1568_),
    .X(_1618_));
 sky130_fd_sc_hd__nand3_1 _2418_ (.A(_1616_),
    .B(_1617_),
    .C(_1568_),
    .Y(_1619_));
 sky130_fd_sc_hd__nand2_1 _2419_ (.A(_1618_),
    .B(_1619_),
    .Y(_1620_));
 sky130_fd_sc_hd__or2_1 _2420_ (.A(_1594_),
    .B(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__nand2_1 _2421_ (.A(_1620_),
    .B(_1594_),
    .Y(_1622_));
 sky130_fd_sc_hd__nand2_2 _2422_ (.A(_1487_),
    .B(_1481_),
    .Y(_1623_));
 sky130_fd_sc_hd__inv_2 _2423_ (.A(_1623_),
    .Y(_1624_));
 sky130_fd_sc_hd__nand2_1 _2424_ (.A(\datapath.MultiplierAC.PPG0.X[4] ),
    .B(_1474_),
    .Y(_1625_));
 sky130_fd_sc_hd__nand2_1 _2425_ (.A(_1624_),
    .B(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__inv_2 _2426_ (.A(_1625_),
    .Y(_1627_));
 sky130_fd_sc_hd__nand2_1 _2427_ (.A(_1627_),
    .B(_1623_),
    .Y(_1628_));
 sky130_fd_sc_hd__nand2_1 _2428_ (.A(_1626_),
    .B(_1628_),
    .Y(_1629_));
 sky130_fd_sc_hd__a21oi_1 _2429_ (.A1(_1572_),
    .A2(_1623_),
    .B1(_1510_),
    .Y(_1630_));
 sky130_fd_sc_hd__nand2_1 _2430_ (.A(_1629_),
    .B(_1630_),
    .Y(_1631_));
 sky130_fd_sc_hd__nand2_1 _2431_ (.A(_1572_),
    .B(_1623_),
    .Y(_1632_));
 sky130_fd_sc_hd__nand2_1 _2432_ (.A(_1632_),
    .B(_1475_),
    .Y(_1633_));
 sky130_fd_sc_hd__nand3_1 _2433_ (.A(_1633_),
    .B(_1626_),
    .C(_1628_),
    .Y(_1634_));
 sky130_fd_sc_hd__nand2_1 _2434_ (.A(_1631_),
    .B(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__inv_2 _2435_ (.A(_1485_),
    .Y(_1636_));
 sky130_fd_sc_hd__nand2_1 _2436_ (.A(_1635_),
    .B(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__nand3_2 _2437_ (.A(_1631_),
    .B(_1634_),
    .C(_1485_),
    .Y(_1638_));
 sky130_fd_sc_hd__nand2_1 _2438_ (.A(_1637_),
    .B(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__inv_2 _2439_ (.A(_1639_),
    .Y(_1640_));
 sky130_fd_sc_hd__nand2_1 _2440_ (.A(_1587_),
    .B(_1583_),
    .Y(_1641_));
 sky130_fd_sc_hd__nand2_1 _2441_ (.A(_1640_),
    .B(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__a21boi_1 _2442_ (.A1(_1580_),
    .A2(_1585_),
    .B1_N(_1583_),
    .Y(_1643_));
 sky130_fd_sc_hd__nand2_1 _2443_ (.A(_1643_),
    .B(_1639_),
    .Y(_1644_));
 sky130_fd_sc_hd__nand2_1 _2444_ (.A(_1642_),
    .B(_1644_),
    .Y(_1645_));
 sky130_fd_sc_hd__nand2_1 _2445_ (.A(_1645_),
    .B(_1623_),
    .Y(_1646_));
 sky130_fd_sc_hd__nand3_1 _2446_ (.A(_1642_),
    .B(_1644_),
    .C(_1624_),
    .Y(_1647_));
 sky130_fd_sc_hd__inv_2 _2447_ (.A(_1589_),
    .Y(_1648_));
 sky130_fd_sc_hd__a21o_1 _2448_ (.A1(_1646_),
    .A2(_1647_),
    .B1(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__nand3_1 _2449_ (.A(_1646_),
    .B(_1647_),
    .C(_1648_),
    .Y(_1650_));
 sky130_fd_sc_hd__a21o_1 _2450_ (.A1(_1649_),
    .A2(_1650_),
    .B1(_1627_),
    .X(_1651_));
 sky130_fd_sc_hd__nand3_1 _2451_ (.A(_1649_),
    .B(_1627_),
    .C(_1650_),
    .Y(_1652_));
 sky130_fd_sc_hd__and3_1 _2452_ (.A(_1651_),
    .B(_1538_),
    .C(_1652_),
    .X(_1653_));
 sky130_fd_sc_hd__a31o_1 _2453_ (.A1(_1621_),
    .A2(_1513_),
    .A3(_1622_),
    .B1(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__nand2_1 _2454_ (.A(_1654_),
    .B(_1517_),
    .Y(_1655_));
 sky130_fd_sc_hd__nand2_1 _2455_ (.A(_1518_),
    .B(_1488_),
    .Y(_1656_));
 sky130_fd_sc_hd__a21oi_1 _2456_ (.A1(_1655_),
    .A2(_1656_),
    .B1(_1545_),
    .Y(_0020_));
 sky130_fd_sc_hd__clkinv_2 _2457_ (.A(_1490_),
    .Y(_1657_));
 sky130_fd_sc_hd__nand2_1 _2458_ (.A(_1613_),
    .B(_1605_),
    .Y(_1658_));
 sky130_fd_sc_hd__nand3_1 _2459_ (.A(_1558_),
    .B(_1547_),
    .C(_1598_),
    .Y(_1659_));
 sky130_fd_sc_hd__a21o_1 _2460_ (.A1(_1527_),
    .A2(_1597_),
    .B1(_1549_),
    .X(_1660_));
 sky130_fd_sc_hd__nand2_1 _2461_ (.A(_1659_),
    .B(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__nand2_1 _2462_ (.A(_1463_),
    .B(\datapath.MultiplierAC.PPG0.X[5] ),
    .Y(_1662_));
 sky130_fd_sc_hd__or2_1 _2463_ (.A(_1597_),
    .B(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__buf_6 _2464_ (.A(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__nand2_1 _2465_ (.A(_1466_),
    .B(\datapath.MultiplierAC.PPG0.X[5] ),
    .Y(_1665_));
 sky130_fd_sc_hd__nand2_1 _2466_ (.A(_1596_),
    .B(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__nand2_1 _2467_ (.A(_1664_),
    .B(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__inv_2 _2468_ (.A(_1667_),
    .Y(_1668_));
 sky130_fd_sc_hd__nand2_1 _2469_ (.A(_1661_),
    .B(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__nand3_1 _2470_ (.A(_1659_),
    .B(_1667_),
    .C(_1660_),
    .Y(_1670_));
 sky130_fd_sc_hd__nand2_1 _2471_ (.A(_1669_),
    .B(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__nand2_1 _2472_ (.A(_1448_),
    .B(_1488_),
    .Y(_1672_));
 sky130_fd_sc_hd__inv_2 _2473_ (.A(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__nand2_1 _2474_ (.A(_1671_),
    .B(_1673_),
    .Y(_1674_));
 sky130_fd_sc_hd__nand3_1 _2475_ (.A(_1669_),
    .B(_1670_),
    .C(_1672_),
    .Y(_1675_));
 sky130_fd_sc_hd__nand2_1 _2476_ (.A(_1674_),
    .B(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__nand2_1 _2477_ (.A(_1658_),
    .B(_1676_),
    .Y(_1677_));
 sky130_fd_sc_hd__nand3b_1 _2478_ (.A_N(_1676_),
    .B(_1613_),
    .C(_1605_),
    .Y(_1678_));
 sky130_fd_sc_hd__nand2_1 _2479_ (.A(_1677_),
    .B(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__nand2_1 _2480_ (.A(_1435_),
    .B(_1485_),
    .Y(_1680_));
 sky130_fd_sc_hd__nand2_1 _2481_ (.A(_1679_),
    .B(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__nand3b_2 _2482_ (.A_N(_1680_),
    .B(_1677_),
    .C(_1678_),
    .Y(_1682_));
 sky130_fd_sc_hd__nand2_1 _2483_ (.A(_1681_),
    .B(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__nand3_1 _2484_ (.A(_1683_),
    .B(_1617_),
    .C(_1619_),
    .Y(_1684_));
 sky130_fd_sc_hd__inv_2 _2485_ (.A(_1683_),
    .Y(_1685_));
 sky130_fd_sc_hd__nand2_1 _2486_ (.A(_1619_),
    .B(_1617_),
    .Y(_1686_));
 sky130_fd_sc_hd__nand2_1 _2487_ (.A(_1685_),
    .B(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__a22o_1 _2488_ (.A1(_1379_),
    .A2(_1475_),
    .B1(_1411_),
    .B2(_1482_),
    .X(_1688_));
 sky130_fd_sc_hd__nand2_1 _2489_ (.A(_1379_),
    .B(_1481_),
    .Y(_1689_));
 sky130_fd_sc_hd__nor2_1 _2490_ (.A(_1594_),
    .B(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__inv_2 _2491_ (.A(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__nand2_1 _2492_ (.A(_1688_),
    .B(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__inv_2 _2493_ (.A(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__a21o_1 _2494_ (.A1(_1684_),
    .A2(_1687_),
    .B1(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__nand3_1 _2495_ (.A(_1684_),
    .B(_1687_),
    .C(_1693_),
    .Y(_1695_));
 sky130_fd_sc_hd__nand2_1 _2496_ (.A(_1694_),
    .B(_1695_),
    .Y(_1696_));
 sky130_fd_sc_hd__or2_1 _2497_ (.A(_1621_),
    .B(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__nand2_1 _2498_ (.A(_1696_),
    .B(_1621_),
    .Y(_1698_));
 sky130_fd_sc_hd__nand3_1 _2499_ (.A(_1697_),
    .B(_1513_),
    .C(_1698_),
    .Y(_1699_));
 sky130_fd_sc_hd__nand2_1 _2500_ (.A(_1650_),
    .B(_1647_),
    .Y(_1700_));
 sky130_fd_sc_hd__nand2_1 _2501_ (.A(_1642_),
    .B(_1638_),
    .Y(_1701_));
 sky130_fd_sc_hd__nand2_1 _2502_ (.A(_1625_),
    .B(_1623_),
    .Y(_1702_));
 sky130_fd_sc_hd__inv_2 _2503_ (.A(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__nand2_1 _2504_ (.A(_1490_),
    .B(_1487_),
    .Y(_1704_));
 sky130_fd_sc_hd__inv_2 _2505_ (.A(_1704_),
    .Y(_1705_));
 sky130_fd_sc_hd__nand2_1 _2506_ (.A(_1575_),
    .B(_1705_),
    .Y(_1706_));
 sky130_fd_sc_hd__o21ai_1 _2507_ (.A1(_1703_),
    .A2(_1633_),
    .B1(_1706_),
    .Y(_1707_));
 sky130_fd_sc_hd__nand2_1 _2508_ (.A(\datapath.MultiplierAC.PPG0.X[5] ),
    .B(\datapath.MultiplierAC.PPG0.X[4] ),
    .Y(_1708_));
 sky130_fd_sc_hd__inv_2 _2509_ (.A(_1708_),
    .Y(_1709_));
 sky130_fd_sc_hd__nand2_1 _2510_ (.A(_1575_),
    .B(_1709_),
    .Y(_1710_));
 sky130_fd_sc_hd__nand2_1 _2511_ (.A(_1492_),
    .B(_1474_),
    .Y(_1711_));
 sky130_fd_sc_hd__nand2_1 _2512_ (.A(_1490_),
    .B(_1481_),
    .Y(_1712_));
 sky130_fd_sc_hd__nand2_1 _2513_ (.A(_1711_),
    .B(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__nand2_1 _2514_ (.A(_1710_),
    .B(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__inv_2 _2515_ (.A(_1714_),
    .Y(_1715_));
 sky130_fd_sc_hd__nand2_1 _2516_ (.A(_1707_),
    .B(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__nand3_1 _2517_ (.A(_1631_),
    .B(_1706_),
    .C(_1714_),
    .Y(_1717_));
 sky130_fd_sc_hd__nand2_1 _2518_ (.A(_1716_),
    .B(_1717_),
    .Y(_1718_));
 sky130_fd_sc_hd__inv_2 _2519_ (.A(_1576_),
    .Y(_1719_));
 sky130_fd_sc_hd__nand2_1 _2520_ (.A(_1718_),
    .B(_1719_),
    .Y(_1720_));
 sky130_fd_sc_hd__nand3_1 _2521_ (.A(_1716_),
    .B(_1717_),
    .C(_1576_),
    .Y(_1721_));
 sky130_fd_sc_hd__nand2_1 _2522_ (.A(_1720_),
    .B(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__nand2_1 _2523_ (.A(_1701_),
    .B(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__nand2_1 _2524_ (.A(_1718_),
    .B(_1576_),
    .Y(_1724_));
 sky130_fd_sc_hd__nand3_1 _2525_ (.A(_1716_),
    .B(_1717_),
    .C(_1719_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_1 _2526_ (.A(_1724_),
    .B(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hd__nand3_1 _2527_ (.A(_1726_),
    .B(_1642_),
    .C(_1638_),
    .Y(_1727_));
 sky130_fd_sc_hd__nand3_2 _2528_ (.A(_1723_),
    .B(_1727_),
    .C(_1719_),
    .Y(_1728_));
 sky130_fd_sc_hd__nand2_1 _2529_ (.A(_1723_),
    .B(_1727_),
    .Y(_1729_));
 sky130_fd_sc_hd__nand2_1 _2530_ (.A(_1729_),
    .B(_1576_),
    .Y(_1730_));
 sky130_fd_sc_hd__nand3_1 _2531_ (.A(_1700_),
    .B(_1728_),
    .C(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__nand2_1 _2532_ (.A(_1730_),
    .B(_1728_),
    .Y(_1732_));
 sky130_fd_sc_hd__a21boi_1 _2533_ (.A1(_1646_),
    .A2(_1648_),
    .B1_N(_1647_),
    .Y(_1733_));
 sky130_fd_sc_hd__nand2_1 _2534_ (.A(_1732_),
    .B(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _2535_ (.A(_1731_),
    .B(_1734_),
    .Y(_1735_));
 sky130_fd_sc_hd__nand2_1 _2536_ (.A(_1735_),
    .B(_1714_),
    .Y(_1736_));
 sky130_fd_sc_hd__nand3_1 _2537_ (.A(_1731_),
    .B(_1734_),
    .C(_1715_),
    .Y(_1737_));
 sky130_fd_sc_hd__nand2_1 _2538_ (.A(_1736_),
    .B(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__or2_1 _2539_ (.A(_1652_),
    .B(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__nand2_1 _2540_ (.A(_1738_),
    .B(_1652_),
    .Y(_1740_));
 sky130_fd_sc_hd__a31oi_1 _2541_ (.A1(_1739_),
    .A2(_1538_),
    .A3(_1740_),
    .B1(_1518_),
    .Y(_1741_));
 sky130_fd_sc_hd__a221oi_1 _2542_ (.A1(_1518_),
    .A2(_1657_),
    .B1(_1699_),
    .B2(_1741_),
    .C1(_1544_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _2543_ (.A(_1652_),
    .Y(_1742_));
 sky130_fd_sc_hd__a21boi_1 _2544_ (.A1(_1736_),
    .A2(_1742_),
    .B1_N(_1737_),
    .Y(_1743_));
 sky130_fd_sc_hd__nand2_1 _2545_ (.A(_1494_),
    .B(_1474_),
    .Y(_1744_));
 sky130_fd_sc_hd__nand2_1 _2546_ (.A(_1582_),
    .B(_1709_),
    .Y(_1745_));
 sky130_fd_sc_hd__nand2_1 _2547_ (.A(_1492_),
    .B(_1481_),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2_1 _2548_ (.A(_1490_),
    .B(_1485_),
    .Y(_1747_));
 sky130_fd_sc_hd__nand2_1 _2549_ (.A(_1746_),
    .B(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__nor2_1 _2550_ (.A(_1574_),
    .B(_1708_),
    .Y(_1749_));
 sky130_fd_sc_hd__a21o_1 _2551_ (.A1(_1745_),
    .A2(_1748_),
    .B1(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__nand3_1 _2552_ (.A(_1745_),
    .B(_1749_),
    .C(_1748_),
    .Y(_1751_));
 sky130_fd_sc_hd__nand2_1 _2553_ (.A(_1750_),
    .B(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__or2_1 _2554_ (.A(_1744_),
    .B(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__nand2_1 _2555_ (.A(_1752_),
    .B(_1744_),
    .Y(_1754_));
 sky130_fd_sc_hd__nand2_1 _2556_ (.A(_1753_),
    .B(_1754_),
    .Y(_1755_));
 sky130_fd_sc_hd__inv_2 _2557_ (.A(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__nand2_1 _2558_ (.A(_1731_),
    .B(_1728_),
    .Y(_1757_));
 sky130_fd_sc_hd__nand3_1 _2559_ (.A(_1722_),
    .B(_1640_),
    .C(_1641_),
    .Y(_1758_));
 sky130_fd_sc_hd__inv_2 _2560_ (.A(_1638_),
    .Y(_1759_));
 sky130_fd_sc_hd__inv_2 _2561_ (.A(_1725_),
    .Y(_1760_));
 sky130_fd_sc_hd__a21oi_1 _2562_ (.A1(_1724_),
    .A2(_1759_),
    .B1(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__nand2_1 _2563_ (.A(_1758_),
    .B(_1761_),
    .Y(_1762_));
 sky130_fd_sc_hd__nand2_1 _2564_ (.A(_1716_),
    .B(_1710_),
    .Y(_1763_));
 sky130_fd_sc_hd__nand2_1 _2565_ (.A(_1494_),
    .B(_1492_),
    .Y(_1764_));
 sky130_fd_sc_hd__nand2_1 _2566_ (.A(_1744_),
    .B(_1746_),
    .Y(_1765_));
 sky130_fd_sc_hd__o21ai_2 _2567_ (.A1(_1574_),
    .A2(_1764_),
    .B1(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hd__inv_2 _2568_ (.A(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__nand2_1 _2569_ (.A(_1763_),
    .B(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__inv_2 _2570_ (.A(_1747_),
    .Y(_1769_));
 sky130_fd_sc_hd__nand3_1 _2571_ (.A(_1716_),
    .B(_1710_),
    .C(_1766_),
    .Y(_1770_));
 sky130_fd_sc_hd__nand3_2 _2572_ (.A(_1768_),
    .B(_1769_),
    .C(_1770_),
    .Y(_1771_));
 sky130_fd_sc_hd__nand2_1 _2573_ (.A(_1763_),
    .B(_1766_),
    .Y(_1772_));
 sky130_fd_sc_hd__nand3_1 _2574_ (.A(_1716_),
    .B(_1710_),
    .C(_1767_),
    .Y(_1773_));
 sky130_fd_sc_hd__nand3_1 _2575_ (.A(_1772_),
    .B(_1747_),
    .C(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__nand2_1 _2576_ (.A(_1771_),
    .B(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__inv_2 _2577_ (.A(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__nand2_1 _2578_ (.A(_1762_),
    .B(_1776_),
    .Y(_1777_));
 sky130_fd_sc_hd__nand3_1 _2579_ (.A(_1775_),
    .B(_1758_),
    .C(_1761_),
    .Y(_1778_));
 sky130_fd_sc_hd__nand2_1 _2580_ (.A(_1777_),
    .B(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__inv_2 _2581_ (.A(_1488_),
    .Y(_1780_));
 sky130_fd_sc_hd__nand2_1 _2582_ (.A(_1779_),
    .B(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hd__nand3_1 _2583_ (.A(_1777_),
    .B(_1778_),
    .C(_1488_),
    .Y(_1782_));
 sky130_fd_sc_hd__nand2_1 _2584_ (.A(_1781_),
    .B(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__nand2_1 _2585_ (.A(_1757_),
    .B(_1783_),
    .Y(_1784_));
 sky130_fd_sc_hd__a21boi_1 _2586_ (.A1(_1700_),
    .A2(_1730_),
    .B1_N(_1728_),
    .Y(_1785_));
 sky130_fd_sc_hd__nand2_1 _2587_ (.A(_1779_),
    .B(_1488_),
    .Y(_1786_));
 sky130_fd_sc_hd__nand3_1 _2588_ (.A(_1777_),
    .B(_1778_),
    .C(_1780_),
    .Y(_1787_));
 sky130_fd_sc_hd__nand2_1 _2589_ (.A(_1786_),
    .B(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hd__nand2_1 _2590_ (.A(_1785_),
    .B(_1788_),
    .Y(_1789_));
 sky130_fd_sc_hd__nand2_1 _2591_ (.A(_1784_),
    .B(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__nor2_1 _2592_ (.A(_1756_),
    .B(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__nand2_1 _2593_ (.A(_1790_),
    .B(_1756_),
    .Y(_1792_));
 sky130_fd_sc_hd__or2b_1 _2594_ (.A(_1791_),
    .B_N(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__or2_1 _2595_ (.A(_1743_),
    .B(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__nand2_1 _2596_ (.A(_1793_),
    .B(_1743_),
    .Y(_1795_));
 sky130_fd_sc_hd__a31o_1 _2597_ (.A1(_1794_),
    .A2(_1538_),
    .A3(_1795_),
    .B1(_1518_),
    .X(_1796_));
 sky130_fd_sc_hd__nand2_1 _2598_ (.A(_1695_),
    .B(_1621_),
    .Y(_1797_));
 sky130_fd_sc_hd__nand2_1 _2599_ (.A(_1694_),
    .B(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__nand2_1 _2600_ (.A(_1687_),
    .B(_1682_),
    .Y(_1799_));
 sky130_fd_sc_hd__nand3_1 _2601_ (.A(_1676_),
    .B(_1611_),
    .C(_1612_),
    .Y(_1800_));
 sky130_fd_sc_hd__nand2_1 _2602_ (.A(_1671_),
    .B(_1672_),
    .Y(_1801_));
 sky130_fd_sc_hd__inv_2 _2603_ (.A(_1605_),
    .Y(_1802_));
 sky130_fd_sc_hd__nand3_1 _2604_ (.A(_1669_),
    .B(_1670_),
    .C(_1673_),
    .Y(_1803_));
 sky130_fd_sc_hd__a21boi_1 _2605_ (.A1(_1801_),
    .A2(_1802_),
    .B1_N(_1803_),
    .Y(_1804_));
 sky130_fd_sc_hd__nand2_1 _2606_ (.A(_1800_),
    .B(_1804_),
    .Y(_1805_));
 sky130_fd_sc_hd__nand2_1 _2607_ (.A(_1669_),
    .B(_1664_),
    .Y(_1806_));
 sky130_fd_sc_hd__nand2_1 _2608_ (.A(_1463_),
    .B(_1494_),
    .Y(_1807_));
 sky130_fd_sc_hd__or2_1 _2609_ (.A(_1665_),
    .B(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__nand2_1 _2610_ (.A(_1466_),
    .B(\datapath.MultiplierAC.PPG0.X[6] ),
    .Y(_1809_));
 sky130_fd_sc_hd__nand2_1 _2611_ (.A(_1662_),
    .B(_1809_),
    .Y(_1810_));
 sky130_fd_sc_hd__nand2_1 _2612_ (.A(_1808_),
    .B(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__inv_2 _2613_ (.A(_1811_),
    .Y(_1812_));
 sky130_fd_sc_hd__nand2_1 _2614_ (.A(_1806_),
    .B(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__nand2_1 _2615_ (.A(_1448_),
    .B(_1490_),
    .Y(_1814_));
 sky130_fd_sc_hd__inv_2 _2616_ (.A(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__nand3_1 _2617_ (.A(_1669_),
    .B(_1664_),
    .C(_1811_),
    .Y(_1816_));
 sky130_fd_sc_hd__nand3_2 _2618_ (.A(_1813_),
    .B(_1815_),
    .C(_1816_),
    .Y(_1817_));
 sky130_fd_sc_hd__nand2_1 _2619_ (.A(_1806_),
    .B(_1811_),
    .Y(_1818_));
 sky130_fd_sc_hd__nand3_1 _2620_ (.A(_1669_),
    .B(_1664_),
    .C(_1812_),
    .Y(_1819_));
 sky130_fd_sc_hd__nand3_1 _2621_ (.A(_1818_),
    .B(_1814_),
    .C(_1819_),
    .Y(_1820_));
 sky130_fd_sc_hd__nand2_1 _2622_ (.A(_1817_),
    .B(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__inv_2 _2623_ (.A(_1821_),
    .Y(_1822_));
 sky130_fd_sc_hd__nand2_1 _2624_ (.A(_1805_),
    .B(_1822_),
    .Y(_1823_));
 sky130_fd_sc_hd__nand3_1 _2625_ (.A(_1821_),
    .B(_1800_),
    .C(_1804_),
    .Y(_1824_));
 sky130_fd_sc_hd__nand2_1 _2626_ (.A(_1823_),
    .B(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__nand2_1 _2627_ (.A(_1435_),
    .B(_1488_),
    .Y(_1826_));
 sky130_fd_sc_hd__inv_2 _2628_ (.A(_1826_),
    .Y(_1827_));
 sky130_fd_sc_hd__nand2_1 _2629_ (.A(_1825_),
    .B(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__nand3_1 _2630_ (.A(_1823_),
    .B(_1824_),
    .C(_1826_),
    .Y(_1829_));
 sky130_fd_sc_hd__nand2_1 _2631_ (.A(_1828_),
    .B(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__nand2_1 _2632_ (.A(_1799_),
    .B(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__inv_2 _2633_ (.A(_1830_),
    .Y(_1832_));
 sky130_fd_sc_hd__nand3_1 _2634_ (.A(_1687_),
    .B(_1832_),
    .C(_1682_),
    .Y(_1833_));
 sky130_fd_sc_hd__nand2_1 _2635_ (.A(_1411_),
    .B(_1484_),
    .Y(_1834_));
 sky130_fd_sc_hd__xnor2_1 _2636_ (.A(_1689_),
    .B(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__or2_1 _2637_ (.A(_1691_),
    .B(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__nand2_1 _2638_ (.A(_1835_),
    .B(_1691_),
    .Y(_1837_));
 sky130_fd_sc_hd__nand2_1 _2639_ (.A(_1836_),
    .B(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__inv_2 _2640_ (.A(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__nand2_1 _2641_ (.A(_1343_),
    .B(_1475_),
    .Y(_1840_));
 sky130_fd_sc_hd__inv_2 _2642_ (.A(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__nand2_1 _2643_ (.A(_1839_),
    .B(_1841_),
    .Y(_1842_));
 sky130_fd_sc_hd__nand2_1 _2644_ (.A(_1838_),
    .B(_1840_),
    .Y(_1843_));
 sky130_fd_sc_hd__nand2_1 _2645_ (.A(_1842_),
    .B(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__a21boi_1 _2646_ (.A1(_1831_),
    .A2(_1833_),
    .B1_N(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__nand2_1 _2647_ (.A(_1831_),
    .B(_1833_),
    .Y(_1846_));
 sky130_fd_sc_hd__or2_1 _2648_ (.A(_1844_),
    .B(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__or2b_1 _2649_ (.A(_1845_),
    .B_N(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__or2_1 _2650_ (.A(_1798_),
    .B(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__nand2_1 _2651_ (.A(_1848_),
    .B(_1798_),
    .Y(_1850_));
 sky130_fd_sc_hd__and3_1 _2652_ (.A(_1849_),
    .B(_1513_),
    .C(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__o221a_1 _2653_ (.A1(_1517_),
    .A2(_1492_),
    .B1(_1796_),
    .B2(_1851_),
    .C1(_1078_),
    .X(_0022_));
 sky130_fd_sc_hd__nand3_1 _2654_ (.A(_1830_),
    .B(_1685_),
    .C(_1686_),
    .Y(_1852_));
 sky130_fd_sc_hd__nand2_1 _2655_ (.A(_1825_),
    .B(_1826_),
    .Y(_1853_));
 sky130_fd_sc_hd__inv_2 _2656_ (.A(_1682_),
    .Y(_1854_));
 sky130_fd_sc_hd__nand3_1 _2657_ (.A(_1823_),
    .B(_1824_),
    .C(_1827_),
    .Y(_1855_));
 sky130_fd_sc_hd__a21boi_1 _2658_ (.A1(_1853_),
    .A2(_1854_),
    .B1_N(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__nand2_1 _2659_ (.A(_1852_),
    .B(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__nand2_1 _2660_ (.A(_1823_),
    .B(_1817_),
    .Y(_1858_));
 sky130_fd_sc_hd__nor2_1 _2661_ (.A(_1667_),
    .B(_1811_),
    .Y(_1859_));
 sky130_fd_sc_hd__nand2_1 _2662_ (.A(_1661_),
    .B(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__nand2_1 _2663_ (.A(_1664_),
    .B(_1808_),
    .Y(_1861_));
 sky130_fd_sc_hd__inv_2 _2664_ (.A(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__nand2_1 _2665_ (.A(_1860_),
    .B(_1862_),
    .Y(_1863_));
 sky130_fd_sc_hd__nand2_1 _2666_ (.A(_1463_),
    .B(_1496_),
    .Y(_1864_));
 sky130_fd_sc_hd__nor2_1 _2667_ (.A(_1809_),
    .B(_1864_),
    .Y(_1865_));
 sky130_fd_sc_hd__clkinv_4 _2668_ (.A(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__nand2_1 _2669_ (.A(_1466_),
    .B(_1496_),
    .Y(_1867_));
 sky130_fd_sc_hd__nand2_1 _2670_ (.A(_1807_),
    .B(_1867_),
    .Y(_1868_));
 sky130_fd_sc_hd__nand2_1 _2671_ (.A(_1866_),
    .B(_1868_),
    .Y(_1869_));
 sky130_fd_sc_hd__inv_2 _2672_ (.A(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__nand2_1 _2673_ (.A(_1863_),
    .B(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__nand3_1 _2674_ (.A(_1860_),
    .B(_1862_),
    .C(_1869_),
    .Y(_1872_));
 sky130_fd_sc_hd__nand2_1 _2675_ (.A(_1871_),
    .B(_1872_),
    .Y(_1873_));
 sky130_fd_sc_hd__nand2_1 _2676_ (.A(_1448_),
    .B(_1492_),
    .Y(_1874_));
 sky130_fd_sc_hd__inv_2 _2677_ (.A(_1874_),
    .Y(_1875_));
 sky130_fd_sc_hd__nand2_1 _2678_ (.A(_1873_),
    .B(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__nand3_1 _2679_ (.A(_1871_),
    .B(_1872_),
    .C(_1874_),
    .Y(_1877_));
 sky130_fd_sc_hd__nand2_1 _2680_ (.A(_1876_),
    .B(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__inv_2 _2681_ (.A(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hd__nand2_1 _2682_ (.A(_1858_),
    .B(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__nand3_1 _2683_ (.A(_1823_),
    .B(_1817_),
    .C(_1878_),
    .Y(_1881_));
 sky130_fd_sc_hd__nand2_1 _2684_ (.A(_1435_),
    .B(_1490_),
    .Y(_1882_));
 sky130_fd_sc_hd__nand3_1 _2685_ (.A(_1880_),
    .B(_1881_),
    .C(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__nand2_1 _2686_ (.A(_1858_),
    .B(_1878_),
    .Y(_1884_));
 sky130_fd_sc_hd__inv_2 _2687_ (.A(_1882_),
    .Y(_1885_));
 sky130_fd_sc_hd__nand3_1 _2688_ (.A(_1823_),
    .B(_1817_),
    .C(_1879_),
    .Y(_1886_));
 sky130_fd_sc_hd__nand3_2 _2689_ (.A(_1884_),
    .B(_1885_),
    .C(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__nand2_1 _2690_ (.A(_1883_),
    .B(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hd__inv_2 _2691_ (.A(_1888_),
    .Y(_1889_));
 sky130_fd_sc_hd__nand2_1 _2692_ (.A(_1857_),
    .B(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__nand3_1 _2693_ (.A(_1852_),
    .B(_1888_),
    .C(_1856_),
    .Y(_1891_));
 sky130_fd_sc_hd__nand2_1 _2694_ (.A(_1890_),
    .B(_1891_),
    .Y(_1892_));
 sky130_fd_sc_hd__nand2_1 _2695_ (.A(_1343_),
    .B(_1482_),
    .Y(_1893_));
 sky130_fd_sc_hd__a22o_1 _2696_ (.A1(_1379_),
    .A2(_1484_),
    .B1(_1411_),
    .B2(_1487_),
    .X(_1894_));
 sky130_fd_sc_hd__nand2_1 _2697_ (.A(_1379_),
    .B(_1487_),
    .Y(_1895_));
 sky130_fd_sc_hd__nor2_1 _2698_ (.A(_1834_),
    .B(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__inv_2 _2699_ (.A(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__a21o_1 _2700_ (.A1(_1594_),
    .A2(_1834_),
    .B1(_1689_),
    .X(_1898_));
 sky130_fd_sc_hd__inv_2 _2701_ (.A(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__a21o_1 _2702_ (.A1(_1894_),
    .A2(_1897_),
    .B1(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__and2_1 _2703_ (.A(_1894_),
    .B(_1897_),
    .X(_1901_));
 sky130_fd_sc_hd__nand2_1 _2704_ (.A(_1901_),
    .B(_1899_),
    .Y(_1902_));
 sky130_fd_sc_hd__nand2_1 _2705_ (.A(_1900_),
    .B(_1902_),
    .Y(_1903_));
 sky130_fd_sc_hd__or2_1 _2706_ (.A(_1893_),
    .B(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__nand2_1 _2707_ (.A(_1903_),
    .B(_1893_),
    .Y(_1905_));
 sky130_fd_sc_hd__nand2_1 _2708_ (.A(_1904_),
    .B(_1905_),
    .Y(_1906_));
 sky130_fd_sc_hd__nand2_1 _2709_ (.A(_1906_),
    .B(_1842_),
    .Y(_1907_));
 sky130_fd_sc_hd__inv_2 _2710_ (.A(_1842_),
    .Y(_1908_));
 sky130_fd_sc_hd__nand3_1 _2711_ (.A(_1904_),
    .B(_1905_),
    .C(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__nand2_1 _2712_ (.A(_1907_),
    .B(_1909_),
    .Y(_1910_));
 sky130_fd_sc_hd__inv_2 _2713_ (.A(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__nand2_1 _2714_ (.A(_1311_),
    .B(_1475_),
    .Y(_1912_));
 sky130_fd_sc_hd__inv_2 _2715_ (.A(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__nand2_1 _2716_ (.A(_1911_),
    .B(_1913_),
    .Y(_1914_));
 sky130_fd_sc_hd__nand2_1 _2717_ (.A(_1910_),
    .B(_1912_),
    .Y(_1915_));
 sky130_fd_sc_hd__nand2_1 _2718_ (.A(_1914_),
    .B(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__nand2_1 _2719_ (.A(_1892_),
    .B(_1916_),
    .Y(_1917_));
 sky130_fd_sc_hd__nand3b_1 _2720_ (.A_N(_1916_),
    .B(_1890_),
    .C(_1891_),
    .Y(_1918_));
 sky130_fd_sc_hd__nand2_1 _2721_ (.A(_1917_),
    .B(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__inv_2 _2722_ (.A(_1919_),
    .Y(_1920_));
 sky130_fd_sc_hd__o21ai_1 _2723_ (.A1(_1798_),
    .A2(_1845_),
    .B1(_1847_),
    .Y(_1921_));
 sky130_fd_sc_hd__or2_1 _2724_ (.A(_1920_),
    .B(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__nand2_1 _2725_ (.A(_1921_),
    .B(_1920_),
    .Y(_1923_));
 sky130_fd_sc_hd__nand2_1 _2726_ (.A(_1777_),
    .B(_1771_),
    .Y(_1924_));
 sky130_fd_sc_hd__nor2_1 _2727_ (.A(_1714_),
    .B(_1766_),
    .Y(_1925_));
 sky130_fd_sc_hd__nand2_1 _2728_ (.A(_1707_),
    .B(_1925_),
    .Y(_1926_));
 sky130_fd_sc_hd__a2bb2oi_1 _2729_ (.A1_N(_1574_),
    .A2_N(_1764_),
    .B1(_1765_),
    .B2(_1749_),
    .Y(_1927_));
 sky130_fd_sc_hd__nand2_1 _2730_ (.A(_1926_),
    .B(_1927_),
    .Y(_1928_));
 sky130_fd_sc_hd__nand2_2 _2731_ (.A(\datapath.MultiplierAC.PPG0.X[7] ),
    .B(\datapath.MultiplierAC.PPG0.X[6] ),
    .Y(_1929_));
 sky130_fd_sc_hd__inv_2 _2732_ (.A(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__nand2_1 _2733_ (.A(_1575_),
    .B(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__nand2_1 _2734_ (.A(\datapath.MultiplierAC.PPG0.X[6] ),
    .B(_1481_),
    .Y(_1932_));
 sky130_fd_sc_hd__nand2_1 _2735_ (.A(_1496_),
    .B(_1474_),
    .Y(_1933_));
 sky130_fd_sc_hd__nand2_1 _2736_ (.A(_1932_),
    .B(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hd__nand2_1 _2737_ (.A(_1931_),
    .B(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__inv_2 _2738_ (.A(_1935_),
    .Y(_1936_));
 sky130_fd_sc_hd__nand2_1 _2739_ (.A(_1928_),
    .B(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__nand3_1 _2740_ (.A(_1926_),
    .B(_1927_),
    .C(_1935_),
    .Y(_1938_));
 sky130_fd_sc_hd__nand2_1 _2741_ (.A(_1937_),
    .B(_1938_),
    .Y(_1939_));
 sky130_fd_sc_hd__nand2_1 _2742_ (.A(_1492_),
    .B(_1485_),
    .Y(_1940_));
 sky130_fd_sc_hd__nand2_1 _2743_ (.A(_1939_),
    .B(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__nand3b_1 _2744_ (.A_N(_1940_),
    .B(_1937_),
    .C(_1938_),
    .Y(_1942_));
 sky130_fd_sc_hd__nand2_1 _2745_ (.A(_1941_),
    .B(_1942_),
    .Y(_1943_));
 sky130_fd_sc_hd__inv_2 _2746_ (.A(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__nand2_1 _2747_ (.A(_1924_),
    .B(_1944_),
    .Y(_1945_));
 sky130_fd_sc_hd__nand3_1 _2748_ (.A(_1777_),
    .B(_1771_),
    .C(_1943_),
    .Y(_1946_));
 sky130_fd_sc_hd__nand2_1 _2749_ (.A(_1945_),
    .B(_1946_),
    .Y(_1947_));
 sky130_fd_sc_hd__nand2_1 _2750_ (.A(_1947_),
    .B(_1704_),
    .Y(_1948_));
 sky130_fd_sc_hd__nand3_1 _2751_ (.A(_1945_),
    .B(_1705_),
    .C(_1946_),
    .Y(_1949_));
 sky130_fd_sc_hd__nand2_1 _2752_ (.A(_1948_),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__nor2_1 _2753_ (.A(_1733_),
    .B(_1732_),
    .Y(_1951_));
 sky130_fd_sc_hd__nand2_1 _2754_ (.A(_1782_),
    .B(_1728_),
    .Y(_1952_));
 sky130_fd_sc_hd__nor2_1 _2755_ (.A(_1951_),
    .B(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__nand2_1 _2756_ (.A(_1950_),
    .B(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__nand3_1 _2757_ (.A(_1731_),
    .B(_1728_),
    .C(_1782_),
    .Y(_1955_));
 sky130_fd_sc_hd__nand3_1 _2758_ (.A(_1955_),
    .B(_1948_),
    .C(_1949_),
    .Y(_1956_));
 sky130_fd_sc_hd__nand2_1 _2759_ (.A(_1954_),
    .B(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__nand2_1 _2760_ (.A(_1719_),
    .B(_1709_),
    .Y(_1958_));
 sky130_fd_sc_hd__nand2_1 _2761_ (.A(_1704_),
    .B(_1940_),
    .Y(_1959_));
 sky130_fd_sc_hd__nand2_1 _2762_ (.A(_1958_),
    .B(_1959_),
    .Y(_1960_));
 sky130_fd_sc_hd__a21o_1 _2763_ (.A1(_1751_),
    .A2(_1745_),
    .B1(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__nand3_1 _2764_ (.A(_1751_),
    .B(_1745_),
    .C(_1960_),
    .Y(_1962_));
 sky130_fd_sc_hd__nand3b_1 _2765_ (.A_N(_1932_),
    .B(_1961_),
    .C(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__nand2_1 _2766_ (.A(_1961_),
    .B(_1962_),
    .Y(_1964_));
 sky130_fd_sc_hd__nand2_1 _2767_ (.A(_1964_),
    .B(_1932_),
    .Y(_1965_));
 sky130_fd_sc_hd__nand3b_1 _2768_ (.A_N(_1753_),
    .B(_1963_),
    .C(_1965_),
    .Y(_1966_));
 sky130_fd_sc_hd__nand2_1 _2769_ (.A(_1965_),
    .B(_1963_),
    .Y(_1967_));
 sky130_fd_sc_hd__nand2_1 _2770_ (.A(_1967_),
    .B(_1753_),
    .Y(_1968_));
 sky130_fd_sc_hd__nand2_1 _2771_ (.A(_1966_),
    .B(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__or2_1 _2772_ (.A(_1933_),
    .B(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__nand2_1 _2773_ (.A(_1969_),
    .B(_1933_),
    .Y(_1971_));
 sky130_fd_sc_hd__nand2_1 _2774_ (.A(_1970_),
    .B(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__inv_2 _2775_ (.A(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__nand2_1 _2776_ (.A(_1957_),
    .B(_1973_),
    .Y(_1974_));
 sky130_fd_sc_hd__nand3_1 _2777_ (.A(_1954_),
    .B(_1956_),
    .C(_1972_),
    .Y(_1975_));
 sky130_fd_sc_hd__nand2_1 _2778_ (.A(_1974_),
    .B(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__o21ai_1 _2779_ (.A1(_1791_),
    .A2(_1743_),
    .B1(_1792_),
    .Y(_1977_));
 sky130_fd_sc_hd__nor2_1 _2780_ (.A(_1976_),
    .B(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__nand2_1 _2781_ (.A(_1977_),
    .B(_1976_),
    .Y(_1979_));
 sky130_fd_sc_hd__and3b_1 _2782_ (.A_N(_1978_),
    .B(_1538_),
    .C(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__a31o_1 _2783_ (.A1(_1513_),
    .A2(_1922_),
    .A3(_1923_),
    .B1(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__nand2_1 _2784_ (.A(_1981_),
    .B(_1517_),
    .Y(_1982_));
 sky130_fd_sc_hd__nand2_1 _2785_ (.A(_1518_),
    .B(_1494_),
    .Y(_1983_));
 sky130_fd_sc_hd__a21oi_1 _2786_ (.A1(_1982_),
    .A2(_1983_),
    .B1(_1545_),
    .Y(_0023_));
 sky130_fd_sc_hd__nand2_1 _2787_ (.A(_1890_),
    .B(_1887_),
    .Y(_1984_));
 sky130_fd_sc_hd__nand3_1 _2788_ (.A(_1805_),
    .B(_1822_),
    .C(_1878_),
    .Y(_1985_));
 sky130_fd_sc_hd__inv_2 _2789_ (.A(_1817_),
    .Y(_1986_));
 sky130_fd_sc_hd__nand2_1 _2790_ (.A(_1873_),
    .B(_1874_),
    .Y(_1987_));
 sky130_fd_sc_hd__nand2_1 _2791_ (.A(_1986_),
    .B(_1987_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2b_1 _2792_ (.A_N(_1873_),
    .B(_1875_),
    .Y(_1989_));
 sky130_fd_sc_hd__and2_1 _2793_ (.A(_1988_),
    .B(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__nand2_1 _2794_ (.A(_1985_),
    .B(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__nand2_1 _2795_ (.A(_1466_),
    .B(_1498_),
    .Y(_1992_));
 sky130_fd_sc_hd__xnor2_1 _2796_ (.A(_1864_),
    .B(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__nor2_1 _2797_ (.A(_1869_),
    .B(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__a2bb2oi_1 _2798_ (.A1_N(_1866_),
    .A2_N(_1993_),
    .B1(_1994_),
    .B2(_1863_),
    .Y(_1995_));
 sky130_fd_sc_hd__nand3_1 _2799_ (.A(_1871_),
    .B(_1866_),
    .C(_1993_),
    .Y(_1996_));
 sky130_fd_sc_hd__nand2_1 _2800_ (.A(_1995_),
    .B(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__nand2_1 _2801_ (.A(_1448_),
    .B(_1494_),
    .Y(_1998_));
 sky130_fd_sc_hd__nand2_1 _2802_ (.A(_1997_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__inv_2 _2803_ (.A(_1998_),
    .Y(_2000_));
 sky130_fd_sc_hd__nand3_2 _2804_ (.A(_1995_),
    .B(_2000_),
    .C(_1996_),
    .Y(_2001_));
 sky130_fd_sc_hd__nand2_1 _2805_ (.A(_1999_),
    .B(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__inv_2 _2806_ (.A(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__nand2_1 _2807_ (.A(_1991_),
    .B(_2003_),
    .Y(_2004_));
 sky130_fd_sc_hd__nand3_1 _2808_ (.A(_1985_),
    .B(_2002_),
    .C(_1990_),
    .Y(_2005_));
 sky130_fd_sc_hd__nand2_1 _2809_ (.A(_2004_),
    .B(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__nand2_1 _2810_ (.A(_1435_),
    .B(_1492_),
    .Y(_2007_));
 sky130_fd_sc_hd__inv_2 _2811_ (.A(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__nand2_1 _2812_ (.A(_2006_),
    .B(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__nand3_1 _2813_ (.A(_2004_),
    .B(_2005_),
    .C(_2007_),
    .Y(_2010_));
 sky130_fd_sc_hd__nand2_1 _2814_ (.A(_2009_),
    .B(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__nand2_1 _2815_ (.A(_1984_),
    .B(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__nand3b_1 _2816_ (.A_N(_2011_),
    .B(_1890_),
    .C(_1887_),
    .Y(_2013_));
 sky130_fd_sc_hd__nand2_1 _2817_ (.A(_2012_),
    .B(_2013_),
    .Y(_2014_));
 sky130_fd_sc_hd__nand2_1 _2818_ (.A(_1902_),
    .B(_1897_),
    .Y(_2015_));
 sky130_fd_sc_hd__nand2_2 _2819_ (.A(_1411_),
    .B(\datapath.MultiplierAC.PPG0.X[4] ),
    .Y(_2016_));
 sky130_fd_sc_hd__xor2_1 _2820_ (.A(_1895_),
    .B(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__nand2_1 _2821_ (.A(_2015_),
    .B(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__nand3b_1 _2822_ (.A_N(_2017_),
    .B(_1902_),
    .C(_1897_),
    .Y(_2019_));
 sky130_fd_sc_hd__nand2_1 _2823_ (.A(_2018_),
    .B(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__inv_2 _2824_ (.A(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__nand2_1 _2825_ (.A(_1343_),
    .B(_1485_),
    .Y(_2022_));
 sky130_fd_sc_hd__inv_2 _2826_ (.A(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__nand2_1 _2827_ (.A(_2021_),
    .B(_2023_),
    .Y(_2024_));
 sky130_fd_sc_hd__nand2_1 _2828_ (.A(_2020_),
    .B(_2022_),
    .Y(_2025_));
 sky130_fd_sc_hd__nand2_1 _2829_ (.A(_2024_),
    .B(_2025_),
    .Y(_2026_));
 sky130_fd_sc_hd__nand3_1 _2830_ (.A(_2026_),
    .B(_1904_),
    .C(_1909_),
    .Y(_2027_));
 sky130_fd_sc_hd__inv_2 _2831_ (.A(_2026_),
    .Y(_2028_));
 sky130_fd_sc_hd__nand2_1 _2832_ (.A(_1909_),
    .B(_1904_),
    .Y(_2029_));
 sky130_fd_sc_hd__nand2_1 _2833_ (.A(_2028_),
    .B(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__nand2_1 _2834_ (.A(_2027_),
    .B(_2030_),
    .Y(_2031_));
 sky130_fd_sc_hd__nand2_1 _2835_ (.A(_1311_),
    .B(_1482_),
    .Y(_2032_));
 sky130_fd_sc_hd__nand2_1 _2836_ (.A(_2031_),
    .B(_2032_),
    .Y(_2033_));
 sky130_fd_sc_hd__nand3b_1 _2837_ (.A_N(_2032_),
    .B(_2027_),
    .C(_2030_),
    .Y(_2034_));
 sky130_fd_sc_hd__nand2_1 _2838_ (.A(_2033_),
    .B(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hd__or2_1 _2839_ (.A(_1914_),
    .B(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__nand2_1 _2840_ (.A(_2035_),
    .B(_1914_),
    .Y(_2037_));
 sky130_fd_sc_hd__nand2_1 _2841_ (.A(_2036_),
    .B(_2037_),
    .Y(_2038_));
 sky130_fd_sc_hd__nand2_1 _2842_ (.A(_2014_),
    .B(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__inv_2 _2843_ (.A(_2038_),
    .Y(_2040_));
 sky130_fd_sc_hd__nand3_2 _2844_ (.A(_2012_),
    .B(_2013_),
    .C(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__nand2_1 _2845_ (.A(_2039_),
    .B(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hd__inv_2 _2846_ (.A(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__nand2_1 _2847_ (.A(_1923_),
    .B(_1918_),
    .Y(_2044_));
 sky130_fd_sc_hd__or2_1 _2848_ (.A(_2043_),
    .B(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__nand2_1 _2849_ (.A(_2044_),
    .B(_2043_),
    .Y(_2046_));
 sky130_fd_sc_hd__nand2_1 _2850_ (.A(\datapath.MultiplierAC.PPG0.Y[8] ),
    .B(_1474_),
    .Y(_2047_));
 sky130_fd_sc_hd__a21bo_1 _2851_ (.A1(_2045_),
    .A2(_2046_),
    .B1_N(_2047_),
    .X(_2048_));
 sky130_fd_sc_hd__nand3b_2 _2852_ (.A_N(_2047_),
    .B(_2045_),
    .C(_2046_),
    .Y(_2049_));
 sky130_fd_sc_hd__nand2_2 _2853_ (.A(_1498_),
    .B(_1474_),
    .Y(_2050_));
 sky130_fd_sc_hd__a21oi_1 _2854_ (.A1(_1945_),
    .A2(_1946_),
    .B1(_1705_),
    .Y(_2051_));
 sky130_fd_sc_hd__o21ai_1 _2855_ (.A1(_1953_),
    .A2(_2051_),
    .B1(_1949_),
    .Y(_2052_));
 sky130_fd_sc_hd__nor2_1 _2856_ (.A(_1775_),
    .B(_1943_),
    .Y(_2053_));
 sky130_fd_sc_hd__nand2_1 _2857_ (.A(_2053_),
    .B(_1762_),
    .Y(_2054_));
 sky130_fd_sc_hd__inv_2 _2858_ (.A(_1771_),
    .Y(_2055_));
 sky130_fd_sc_hd__a21boi_1 _2859_ (.A1(_2055_),
    .A2(_1941_),
    .B1_N(_1942_),
    .Y(_2056_));
 sky130_fd_sc_hd__nand2_1 _2860_ (.A(_2054_),
    .B(_2056_),
    .Y(_2057_));
 sky130_fd_sc_hd__nand2_1 _2861_ (.A(_1937_),
    .B(_1931_),
    .Y(_2058_));
 sky130_fd_sc_hd__nand2_1 _2862_ (.A(_1498_),
    .B(\datapath.MultiplierAC.PPG0.X[7] ),
    .Y(_2059_));
 sky130_fd_sc_hd__inv_2 _2863_ (.A(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__nand2_1 _2864_ (.A(_1575_),
    .B(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__nand2_1 _2865_ (.A(_1496_),
    .B(_1481_),
    .Y(_2062_));
 sky130_fd_sc_hd__nand2_1 _2866_ (.A(_2050_),
    .B(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__nand2_1 _2867_ (.A(_2061_),
    .B(_2063_),
    .Y(_2064_));
 sky130_fd_sc_hd__nand2_1 _2868_ (.A(_2058_),
    .B(_2064_),
    .Y(_2065_));
 sky130_fd_sc_hd__inv_2 _2869_ (.A(_2064_),
    .Y(_2066_));
 sky130_fd_sc_hd__nand3_1 _2870_ (.A(_1937_),
    .B(_1931_),
    .C(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__nand2_1 _2871_ (.A(_2065_),
    .B(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__nand2_1 _2872_ (.A(_1494_),
    .B(_1485_),
    .Y(_2069_));
 sky130_fd_sc_hd__inv_2 _2873_ (.A(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__nand2_1 _2874_ (.A(_2068_),
    .B(_2070_),
    .Y(_2071_));
 sky130_fd_sc_hd__nand3_1 _2875_ (.A(_2065_),
    .B(_2069_),
    .C(_2067_),
    .Y(_2072_));
 sky130_fd_sc_hd__nand2_1 _2876_ (.A(_2071_),
    .B(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__inv_2 _2877_ (.A(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__nand2_1 _2878_ (.A(_2057_),
    .B(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__nand3_1 _2879_ (.A(_2054_),
    .B(_2073_),
    .C(_2056_),
    .Y(_2076_));
 sky130_fd_sc_hd__nand2_1 _2880_ (.A(_2075_),
    .B(_2076_),
    .Y(_2077_));
 sky130_fd_sc_hd__nand2_1 _2881_ (.A(_1492_),
    .B(_1487_),
    .Y(_2078_));
 sky130_fd_sc_hd__nand2_1 _2882_ (.A(_2077_),
    .B(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hd__nand3b_1 _2883_ (.A_N(_2078_),
    .B(_2075_),
    .C(_2076_),
    .Y(_2080_));
 sky130_fd_sc_hd__nand2_1 _2884_ (.A(_2079_),
    .B(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__inv_2 _2885_ (.A(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__nand2_1 _2886_ (.A(_2052_),
    .B(_2082_),
    .Y(_2083_));
 sky130_fd_sc_hd__nand3_1 _2887_ (.A(_1956_),
    .B(_2081_),
    .C(_1949_),
    .Y(_2084_));
 sky130_fd_sc_hd__nand2_1 _2888_ (.A(_2083_),
    .B(_2084_),
    .Y(_2085_));
 sky130_fd_sc_hd__nand2_1 _2889_ (.A(_1961_),
    .B(_1958_),
    .Y(_2086_));
 sky130_fd_sc_hd__nand2_1 _2890_ (.A(_1709_),
    .B(_1488_),
    .Y(_2087_));
 sky130_fd_sc_hd__nand2_1 _2891_ (.A(_2078_),
    .B(_1657_),
    .Y(_2088_));
 sky130_fd_sc_hd__nand2_1 _2892_ (.A(_2087_),
    .B(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__nand2_1 _2893_ (.A(_2086_),
    .B(_2089_),
    .Y(_2090_));
 sky130_fd_sc_hd__inv_2 _2894_ (.A(_2089_),
    .Y(_2091_));
 sky130_fd_sc_hd__nand3_1 _2895_ (.A(_1961_),
    .B(_1958_),
    .C(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__nand2_1 _2896_ (.A(_2090_),
    .B(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__nand2_1 _2897_ (.A(_2093_),
    .B(_2070_),
    .Y(_2094_));
 sky130_fd_sc_hd__nand3_1 _2898_ (.A(_2090_),
    .B(_2069_),
    .C(_2092_),
    .Y(_2095_));
 sky130_fd_sc_hd__nand2_1 _2899_ (.A(_2094_),
    .B(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__nand3_1 _2900_ (.A(_2096_),
    .B(_1963_),
    .C(_1966_),
    .Y(_2097_));
 sky130_fd_sc_hd__inv_2 _2901_ (.A(_2096_),
    .Y(_2098_));
 sky130_fd_sc_hd__nand2_1 _2902_ (.A(_1966_),
    .B(_1963_),
    .Y(_2099_));
 sky130_fd_sc_hd__nand2_1 _2903_ (.A(_2098_),
    .B(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__nand2_1 _2904_ (.A(_2097_),
    .B(_2100_),
    .Y(_2101_));
 sky130_fd_sc_hd__nand2_1 _2905_ (.A(_2101_),
    .B(_2062_),
    .Y(_2102_));
 sky130_fd_sc_hd__nand3b_1 _2906_ (.A_N(_2062_),
    .B(_2097_),
    .C(_2100_),
    .Y(_2103_));
 sky130_fd_sc_hd__nand2_1 _2907_ (.A(_2102_),
    .B(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__or2_1 _2908_ (.A(_1970_),
    .B(_2104_),
    .X(_2105_));
 sky130_fd_sc_hd__nand2_1 _2909_ (.A(_2104_),
    .B(_1970_),
    .Y(_2106_));
 sky130_fd_sc_hd__nand2_1 _2910_ (.A(_2105_),
    .B(_2106_),
    .Y(_2107_));
 sky130_fd_sc_hd__nand2_1 _2911_ (.A(_2085_),
    .B(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__inv_2 _2912_ (.A(_2107_),
    .Y(_2109_));
 sky130_fd_sc_hd__nand3_1 _2913_ (.A(_2083_),
    .B(_2109_),
    .C(_2084_),
    .Y(_2110_));
 sky130_fd_sc_hd__nand2_1 _2914_ (.A(_2108_),
    .B(_2110_),
    .Y(_2111_));
 sky130_fd_sc_hd__inv_2 _2915_ (.A(_2111_),
    .Y(_2112_));
 sky130_fd_sc_hd__or2_1 _2916_ (.A(_1972_),
    .B(_1957_),
    .X(_2113_));
 sky130_fd_sc_hd__nand2_1 _2917_ (.A(_1979_),
    .B(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__or2_1 _2918_ (.A(_2112_),
    .B(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__nand2_1 _2919_ (.A(_2114_),
    .B(_2112_),
    .Y(_2116_));
 sky130_fd_sc_hd__nand2_1 _2920_ (.A(_2115_),
    .B(_2116_),
    .Y(_2117_));
 sky130_fd_sc_hd__nor2_1 _2921_ (.A(_2050_),
    .B(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__inv_2 _2922_ (.A(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__nand2_1 _2923_ (.A(_2117_),
    .B(_2050_),
    .Y(_2120_));
 sky130_fd_sc_hd__and3_1 _2924_ (.A(_2119_),
    .B(_1538_),
    .C(_2120_),
    .X(_2121_));
 sky130_fd_sc_hd__a31o_1 _2925_ (.A1(_2048_),
    .A2(_1513_),
    .A3(_2049_),
    .B1(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__nand2_1 _2926_ (.A(_2122_),
    .B(_1517_),
    .Y(_2123_));
 sky130_fd_sc_hd__nand2_1 _2927_ (.A(_1518_),
    .B(_1496_),
    .Y(_2124_));
 sky130_fd_sc_hd__a21oi_1 _2928_ (.A1(_2123_),
    .A2(_2124_),
    .B1(_1545_),
    .Y(_0024_));
 sky130_fd_sc_hd__a22o_1 _2929_ (.A1(_1500_),
    .A2(_1474_),
    .B1(_1498_),
    .B2(_1482_),
    .X(_2125_));
 sky130_fd_sc_hd__nand2_2 _2930_ (.A(_1500_),
    .B(_1498_),
    .Y(_2126_));
 sky130_fd_sc_hd__nor2_1 _2931_ (.A(_1574_),
    .B(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__inv_2 _2932_ (.A(_2127_),
    .Y(_2128_));
 sky130_fd_sc_hd__nand2_1 _2933_ (.A(_2125_),
    .B(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hd__nand2_1 _2934_ (.A(_2116_),
    .B(_2110_),
    .Y(_2130_));
 sky130_fd_sc_hd__nand2_1 _2935_ (.A(_2083_),
    .B(_2080_),
    .Y(_2131_));
 sky130_fd_sc_hd__nand2_1 _2936_ (.A(_2075_),
    .B(_2071_),
    .Y(_2132_));
 sky130_fd_sc_hd__inv_2 _2937_ (.A(_2129_),
    .Y(_2133_));
 sky130_fd_sc_hd__nand2_1 _2938_ (.A(_1936_),
    .B(_2066_),
    .Y(_2134_));
 sky130_fd_sc_hd__and2_1 _2939_ (.A(_1931_),
    .B(_2061_),
    .X(_2135_));
 sky130_fd_sc_hd__o21a_1 _2940_ (.A1(_2134_),
    .A2(_1927_),
    .B1(_2135_),
    .X(_2136_));
 sky130_fd_sc_hd__nand3b_1 _2941_ (.A_N(_2134_),
    .B(_1707_),
    .C(_1925_),
    .Y(_2137_));
 sky130_fd_sc_hd__nand2_1 _2942_ (.A(_2136_),
    .B(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__or2_1 _2943_ (.A(_2133_),
    .B(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__nand2_1 _2944_ (.A(_2138_),
    .B(_2133_),
    .Y(_2140_));
 sky130_fd_sc_hd__nand2_1 _2945_ (.A(_1496_),
    .B(_1485_),
    .Y(_2141_));
 sky130_fd_sc_hd__inv_2 _2946_ (.A(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__a21o_1 _2947_ (.A1(_2139_),
    .A2(_2140_),
    .B1(_2142_),
    .X(_2143_));
 sky130_fd_sc_hd__nand3_1 _2948_ (.A(_2139_),
    .B(_2142_),
    .C(_2140_),
    .Y(_2144_));
 sky130_fd_sc_hd__nand2_1 _2949_ (.A(_2143_),
    .B(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__inv_2 _2950_ (.A(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__nand2_1 _2951_ (.A(_2132_),
    .B(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__nand3_1 _2952_ (.A(_2145_),
    .B(_2075_),
    .C(_2071_),
    .Y(_2148_));
 sky130_fd_sc_hd__nand2_1 _2953_ (.A(_2147_),
    .B(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__nand2_1 _2954_ (.A(_1494_),
    .B(_1488_),
    .Y(_2150_));
 sky130_fd_sc_hd__nand2_1 _2955_ (.A(_2149_),
    .B(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__inv_2 _2956_ (.A(_2150_),
    .Y(_2152_));
 sky130_fd_sc_hd__nand3_1 _2957_ (.A(_2147_),
    .B(_2148_),
    .C(_2152_),
    .Y(_2153_));
 sky130_fd_sc_hd__nand2_1 _2958_ (.A(_2151_),
    .B(_2153_),
    .Y(_2154_));
 sky130_fd_sc_hd__inv_2 _2959_ (.A(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__nand2_1 _2960_ (.A(_2131_),
    .B(_2155_),
    .Y(_2156_));
 sky130_fd_sc_hd__nand3_1 _2961_ (.A(_2083_),
    .B(_2154_),
    .C(_2080_),
    .Y(_2157_));
 sky130_fd_sc_hd__nand2_1 _2962_ (.A(_2156_),
    .B(_2157_),
    .Y(_2158_));
 sky130_fd_sc_hd__inv_2 _2963_ (.A(_1970_),
    .Y(_2159_));
 sky130_fd_sc_hd__a21boi_1 _2964_ (.A1(_2102_),
    .A2(_2159_),
    .B1_N(_2103_),
    .Y(_2160_));
 sky130_fd_sc_hd__nand2_1 _2965_ (.A(_2100_),
    .B(_2094_),
    .Y(_2161_));
 sky130_fd_sc_hd__nand2_1 _2966_ (.A(_1961_),
    .B(_2087_),
    .Y(_2162_));
 sky130_fd_sc_hd__or2_1 _2967_ (.A(_2152_),
    .B(_2162_),
    .X(_2163_));
 sky130_fd_sc_hd__nand2_1 _2968_ (.A(_2162_),
    .B(_2152_),
    .Y(_2164_));
 sky130_fd_sc_hd__nand2_1 _2969_ (.A(_2163_),
    .B(_2164_),
    .Y(_2165_));
 sky130_fd_sc_hd__inv_2 _2970_ (.A(_2165_),
    .Y(_2166_));
 sky130_fd_sc_hd__nand2_1 _2971_ (.A(_2161_),
    .B(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__nand3_1 _2972_ (.A(_2100_),
    .B(_2094_),
    .C(_2165_),
    .Y(_2168_));
 sky130_fd_sc_hd__nand2_1 _2973_ (.A(_2167_),
    .B(_2168_),
    .Y(_2169_));
 sky130_fd_sc_hd__xor2_1 _2974_ (.A(_2142_),
    .B(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__xor2_1 _2975_ (.A(_2160_),
    .B(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__inv_2 _2976_ (.A(_2171_),
    .Y(_2172_));
 sky130_fd_sc_hd__nand2_1 _2977_ (.A(_2158_),
    .B(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__nand3_1 _2978_ (.A(_2156_),
    .B(_2171_),
    .C(_2157_),
    .Y(_2174_));
 sky130_fd_sc_hd__nand2_1 _2979_ (.A(_2173_),
    .B(_2174_),
    .Y(_2175_));
 sky130_fd_sc_hd__inv_2 _2980_ (.A(_2175_),
    .Y(_2176_));
 sky130_fd_sc_hd__nand2_1 _2981_ (.A(_2130_),
    .B(_2176_),
    .Y(_2177_));
 sky130_fd_sc_hd__nand3_1 _2982_ (.A(_2175_),
    .B(_2116_),
    .C(_2110_),
    .Y(_2178_));
 sky130_fd_sc_hd__nand2_1 _2983_ (.A(_2177_),
    .B(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__nor2_1 _2984_ (.A(_2129_),
    .B(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hd__nand2_1 _2985_ (.A(_2179_),
    .B(_2129_),
    .Y(_2181_));
 sky130_fd_sc_hd__or2b_1 _2986_ (.A(_2180_),
    .B_N(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__nand2_1 _2987_ (.A(_2182_),
    .B(_2119_),
    .Y(_2183_));
 sky130_fd_sc_hd__or2_1 _2988_ (.A(_2119_),
    .B(_2182_),
    .X(_2184_));
 sky130_fd_sc_hd__nand2_1 _2989_ (.A(_2046_),
    .B(_2041_),
    .Y(_2185_));
 sky130_fd_sc_hd__nand3_1 _2990_ (.A(_1857_),
    .B(_2011_),
    .C(_1889_),
    .Y(_2186_));
 sky130_fd_sc_hd__nand2_1 _2991_ (.A(_2006_),
    .B(_2007_),
    .Y(_2187_));
 sky130_fd_sc_hd__inv_2 _2992_ (.A(_1887_),
    .Y(_2188_));
 sky130_fd_sc_hd__nand3_1 _2993_ (.A(_2004_),
    .B(_2005_),
    .C(_2008_),
    .Y(_2189_));
 sky130_fd_sc_hd__a21boi_1 _2994_ (.A1(_2187_),
    .A2(_2188_),
    .B1_N(_2189_),
    .Y(_2190_));
 sky130_fd_sc_hd__nand2_1 _2995_ (.A(_2186_),
    .B(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__nand2_1 _2996_ (.A(_2004_),
    .B(_2001_),
    .Y(_2192_));
 sky130_fd_sc_hd__nand3_1 _2997_ (.A(_1661_),
    .B(_1994_),
    .C(_1859_),
    .Y(_2193_));
 sky130_fd_sc_hd__nand2_1 _2998_ (.A(_1994_),
    .B(_1861_),
    .Y(_0080_));
 sky130_fd_sc_hd__a21o_1 _2999_ (.A1(_1809_),
    .A2(_1992_),
    .B1(_1864_),
    .X(_0081_));
 sky130_fd_sc_hd__nand2_1 _3000_ (.A(_0080_),
    .B(_0081_),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _3001_ (.A(_0082_),
    .Y(_0083_));
 sky130_fd_sc_hd__nand2_1 _3002_ (.A(_2193_),
    .B(_0083_),
    .Y(_0084_));
 sky130_fd_sc_hd__a22o_1 _3003_ (.A1(_1463_),
    .A2(_1498_),
    .B1(_1466_),
    .B2(_1500_),
    .X(_0085_));
 sky130_fd_sc_hd__nand2_1 _3004_ (.A(_1463_),
    .B(_1500_),
    .Y(_0086_));
 sky130_fd_sc_hd__nor2_1 _3005_ (.A(_1992_),
    .B(_0086_),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _3006_ (.A(_0087_),
    .Y(_0088_));
 sky130_fd_sc_hd__nand2_1 _3007_ (.A(_0085_),
    .B(_0088_),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _3008_ (.A(_0089_),
    .Y(_0090_));
 sky130_fd_sc_hd__nand2_1 _3009_ (.A(_0084_),
    .B(_0090_),
    .Y(_0091_));
 sky130_fd_sc_hd__nand3_1 _3010_ (.A(_2193_),
    .B(_0083_),
    .C(_0089_),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_1 _3011_ (.A(_0091_),
    .B(_0092_),
    .Y(_0093_));
 sky130_fd_sc_hd__nand2_1 _3012_ (.A(_1448_),
    .B(_1496_),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _3013_ (.A(_0094_),
    .Y(_0095_));
 sky130_fd_sc_hd__nand2_1 _3014_ (.A(_0093_),
    .B(_0095_),
    .Y(_0096_));
 sky130_fd_sc_hd__nand3_1 _3015_ (.A(_0091_),
    .B(_0092_),
    .C(_0094_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand2_1 _3016_ (.A(_0096_),
    .B(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__nand2_1 _3017_ (.A(_2192_),
    .B(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__nand2_1 _3018_ (.A(_1435_),
    .B(_1494_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _3019_ (.A(_0100_),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _3020_ (.A(_0098_),
    .Y(_0102_));
 sky130_fd_sc_hd__nand3_1 _3021_ (.A(_2004_),
    .B(_2001_),
    .C(_0102_),
    .Y(_0103_));
 sky130_fd_sc_hd__nand3_2 _3022_ (.A(_0099_),
    .B(_0101_),
    .C(_0103_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand2_1 _3023_ (.A(_2192_),
    .B(_0102_),
    .Y(_0105_));
 sky130_fd_sc_hd__nand3_1 _3024_ (.A(_2004_),
    .B(_2001_),
    .C(_0098_),
    .Y(_0106_));
 sky130_fd_sc_hd__nand3_1 _3025_ (.A(_0105_),
    .B(_0100_),
    .C(_0106_),
    .Y(_0107_));
 sky130_fd_sc_hd__nand2_1 _3026_ (.A(_0104_),
    .B(_0107_),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _3027_ (.A(_0108_),
    .Y(_0109_));
 sky130_fd_sc_hd__nand2_1 _3028_ (.A(_2191_),
    .B(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__nand3_1 _3029_ (.A(_2186_),
    .B(_0108_),
    .C(_2190_),
    .Y(_0111_));
 sky130_fd_sc_hd__nand2_1 _3030_ (.A(_0110_),
    .B(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _3031_ (.A(_1914_),
    .Y(_0113_));
 sky130_fd_sc_hd__a21boi_2 _3032_ (.A1(_2033_),
    .A2(_0113_),
    .B1_N(_2034_),
    .Y(_0114_));
 sky130_fd_sc_hd__nand2_1 _3033_ (.A(_1311_),
    .B(_1485_),
    .Y(_0115_));
 sky130_fd_sc_hd__nand2_1 _3034_ (.A(_2030_),
    .B(_2024_),
    .Y(_0116_));
 sky130_fd_sc_hd__nand3_1 _3035_ (.A(_1901_),
    .B(_1899_),
    .C(_2017_),
    .Y(_0117_));
 sky130_fd_sc_hd__a21o_1 _3036_ (.A1(_1834_),
    .A2(_2016_),
    .B1(_1895_),
    .X(_0118_));
 sky130_fd_sc_hd__nand2_1 _3037_ (.A(_0117_),
    .B(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__a22o_1 _3038_ (.A1(_1379_),
    .A2(_1490_),
    .B1(_1411_),
    .B2(_1492_),
    .X(_0120_));
 sky130_fd_sc_hd__nand2_1 _3039_ (.A(_1379_),
    .B(\datapath.MultiplierAC.PPG0.X[5] ),
    .Y(_0121_));
 sky130_fd_sc_hd__nor2_1 _3040_ (.A(_2016_),
    .B(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _3041_ (.A(_0122_),
    .Y(_0123_));
 sky130_fd_sc_hd__nand2_1 _3042_ (.A(_0120_),
    .B(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__nand2b_1 _3043_ (.A_N(_0119_),
    .B(_0124_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _3044_ (.A(_0124_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_1 _3045_ (.A(_0119_),
    .B(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__nand2_1 _3046_ (.A(_0125_),
    .B(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__nand2_1 _3047_ (.A(_1343_),
    .B(_1488_),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _3048_ (.A(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__nand2_1 _3049_ (.A(_0128_),
    .B(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__nand3_1 _3050_ (.A(_0125_),
    .B(_0127_),
    .C(_0129_),
    .Y(_0132_));
 sky130_fd_sc_hd__nand2_1 _3051_ (.A(_0131_),
    .B(_0132_),
    .Y(_0133_));
 sky130_fd_sc_hd__nand2_1 _3052_ (.A(_0116_),
    .B(_0133_),
    .Y(_0134_));
 sky130_fd_sc_hd__nand2_1 _3053_ (.A(_0128_),
    .B(_0129_),
    .Y(_0135_));
 sky130_fd_sc_hd__nand3_1 _3054_ (.A(_0125_),
    .B(_0127_),
    .C(_0130_),
    .Y(_0136_));
 sky130_fd_sc_hd__nand2_1 _3055_ (.A(_0135_),
    .B(_0136_),
    .Y(_0137_));
 sky130_fd_sc_hd__nand3_1 _3056_ (.A(_2030_),
    .B(_2024_),
    .C(_0137_),
    .Y(_0138_));
 sky130_fd_sc_hd__nand2_1 _3057_ (.A(_0134_),
    .B(_0138_),
    .Y(_0139_));
 sky130_fd_sc_hd__nor2_1 _3058_ (.A(_0115_),
    .B(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _3059_ (.A(_0140_),
    .Y(_0141_));
 sky130_fd_sc_hd__nand2_1 _3060_ (.A(_0139_),
    .B(_0115_),
    .Y(_0142_));
 sky130_fd_sc_hd__nand2_1 _3061_ (.A(_0141_),
    .B(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__xor2_2 _3062_ (.A(_0114_),
    .B(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__inv_2 _3063_ (.A(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__nand2_1 _3064_ (.A(_0112_),
    .B(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__nand3_1 _3065_ (.A(_0110_),
    .B(_0144_),
    .C(_0111_),
    .Y(_0147_));
 sky130_fd_sc_hd__nand2_1 _3066_ (.A(_0146_),
    .B(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__nand2_1 _3068_ (.A(_2185_),
    .B(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__nand3_1 _3069_ (.A(_2046_),
    .B(_2041_),
    .C(_0148_),
    .Y(_0151_));
 sky130_fd_sc_hd__nand2_1 _3070_ (.A(_0150_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__a22o_1 _3071_ (.A1(\datapath.MultiplierAC.PPG0.Y[9] ),
    .A2(_1475_),
    .B1(\datapath.MultiplierAC.PPG0.Y[8] ),
    .B2(_1482_),
    .X(_0153_));
 sky130_fd_sc_hd__nand2_1 _3072_ (.A(\datapath.MultiplierAC.PPG0.Y[9] ),
    .B(_1481_),
    .Y(_0154_));
 sky130_fd_sc_hd__nor2_1 _3073_ (.A(_2047_),
    .B(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _3074_ (.A(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__nand2_1 _3075_ (.A(_0153_),
    .B(_0156_),
    .Y(_0157_));
 sky130_fd_sc_hd__nand2_1 _3076_ (.A(_0152_),
    .B(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _3077_ (.A(_0157_),
    .Y(_0159_));
 sky130_fd_sc_hd__nand3_1 _3078_ (.A(_0150_),
    .B(_0151_),
    .C(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__nand2_1 _3079_ (.A(_0158_),
    .B(_0160_),
    .Y(_0161_));
 sky130_fd_sc_hd__xor2_1 _3080_ (.A(_2049_),
    .B(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__a32o_1 _3081_ (.A1(_1538_),
    .A2(_2183_),
    .A3(_2184_),
    .B1(_0162_),
    .B2(_1513_),
    .X(_0163_));
 sky130_fd_sc_hd__nand2_1 _3082_ (.A(_0163_),
    .B(_1517_),
    .Y(_0164_));
 sky130_fd_sc_hd__nand2_1 _3083_ (.A(_1518_),
    .B(_1498_),
    .Y(_0165_));
 sky130_fd_sc_hd__a21oi_1 _3084_ (.A1(_0164_),
    .A2(_0165_),
    .B1(_1545_),
    .Y(_0025_));
 sky130_fd_sc_hd__nand2_1 _3085_ (.A(_0160_),
    .B(_2049_),
    .Y(_0166_));
 sky130_fd_sc_hd__nand2_1 _3086_ (.A(_0166_),
    .B(_0158_),
    .Y(_0167_));
 sky130_fd_sc_hd__nand3_1 _3087_ (.A(_0149_),
    .B(_2043_),
    .C(_2044_),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _3088_ (.A(_2041_),
    .Y(_0169_));
 sky130_fd_sc_hd__a21boi_1 _3089_ (.A1(_0146_),
    .A2(_0169_),
    .B1_N(_0147_),
    .Y(_0170_));
 sky130_fd_sc_hd__nand2_1 _3090_ (.A(_0168_),
    .B(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__nand2_1 _3091_ (.A(_0110_),
    .B(_0104_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand3_1 _3092_ (.A(_1999_),
    .B(_0098_),
    .C(_2001_),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _3093_ (.A(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__nand2_1 _3094_ (.A(_0174_),
    .B(_1991_),
    .Y(_0175_));
 sky130_fd_sc_hd__or2_1 _3095_ (.A(_0094_),
    .B(_0093_),
    .X(_0176_));
 sky130_fd_sc_hd__o21a_1 _3096_ (.A1(_2001_),
    .A2(_0102_),
    .B1(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _3097_ (.A(_0175_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand2_1 _3098_ (.A(_1466_),
    .B(_1502_),
    .Y(_0179_));
 sky130_fd_sc_hd__nor2_1 _3099_ (.A(_0086_),
    .B(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_1 _3100_ (.A(_0086_),
    .B(_0179_),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _3101_ (.A(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__nor2_1 _3102_ (.A(_0180_),
    .B(_0182_),
    .Y(_0183_));
 sky130_fd_sc_hd__nand2_1 _3103_ (.A(_0091_),
    .B(_0088_),
    .Y(_0184_));
 sky130_fd_sc_hd__xor2_1 _3104_ (.A(_0183_),
    .B(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__nand3_1 _3105_ (.A(_0185_),
    .B(_1448_),
    .C(_1498_),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _3106_ (.A(_1498_),
    .Y(_0187_));
 sky130_fd_sc_hd__xnor2_1 _3107_ (.A(_0183_),
    .B(_0184_),
    .Y(_0188_));
 sky130_fd_sc_hd__o21ai_1 _3108_ (.A1(_1457_),
    .A2(_0187_),
    .B1(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__nand2_1 _3109_ (.A(_0186_),
    .B(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _3110_ (.A(_0190_),
    .Y(_0191_));
 sky130_fd_sc_hd__nand2_1 _3111_ (.A(_0178_),
    .B(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__nand3_1 _3112_ (.A(_0190_),
    .B(_0175_),
    .C(_0177_),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2_1 _3113_ (.A(_0192_),
    .B(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__nand2_1 _3114_ (.A(_1435_),
    .B(_1496_),
    .Y(_0195_));
 sky130_fd_sc_hd__nand2_1 _3115_ (.A(_0194_),
    .B(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__nand3b_1 _3116_ (.A_N(_0195_),
    .B(_0192_),
    .C(_0193_),
    .Y(_0197_));
 sky130_fd_sc_hd__nand2_1 _3117_ (.A(_0196_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__nand2_1 _3118_ (.A(_0172_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__inv_2 _3119_ (.A(_0198_),
    .Y(_0200_));
 sky130_fd_sc_hd__nand3_1 _3120_ (.A(_0110_),
    .B(_0104_),
    .C(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__nand2_1 _3121_ (.A(_0199_),
    .B(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__nand3_1 _3122_ (.A(_0133_),
    .B(_2028_),
    .C(_2029_),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_2 _3123_ (.A(_2024_),
    .Y(_0204_));
 sky130_fd_sc_hd__a21boi_1 _3124_ (.A1(_0135_),
    .A2(_0204_),
    .B1_N(_0136_),
    .Y(_0205_));
 sky130_fd_sc_hd__nand2_1 _3125_ (.A(_0203_),
    .B(_0205_),
    .Y(_0206_));
 sky130_fd_sc_hd__nand2_1 _3126_ (.A(_1343_),
    .B(_1490_),
    .Y(_0207_));
 sky130_fd_sc_hd__nand2_1 _3127_ (.A(_1411_),
    .B(_1494_),
    .Y(_0208_));
 sky130_fd_sc_hd__nor2_1 _3128_ (.A(_0121_),
    .B(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_2 _3129_ (.A(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__nand2_1 _3130_ (.A(_0121_),
    .B(_0208_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _3131_ (.A(_0210_),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _3132_ (.A(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__nand2_1 _3133_ (.A(_0127_),
    .B(_0123_),
    .Y(_0214_));
 sky130_fd_sc_hd__or2_1 _3134_ (.A(_0213_),
    .B(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__nand2_1 _3135_ (.A(_0214_),
    .B(_0213_),
    .Y(_0216_));
 sky130_fd_sc_hd__nand3b_2 _3136_ (.A_N(_0207_),
    .B(_0215_),
    .C(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _3137_ (.A(_0215_),
    .B(_0216_),
    .Y(_0218_));
 sky130_fd_sc_hd__nand2_1 _3138_ (.A(_0218_),
    .B(_0207_),
    .Y(_0219_));
 sky130_fd_sc_hd__nand3_2 _3139_ (.A(_0206_),
    .B(_0217_),
    .C(_0219_),
    .Y(_0220_));
 sky130_fd_sc_hd__nand2_1 _3140_ (.A(_0219_),
    .B(_0217_),
    .Y(_0221_));
 sky130_fd_sc_hd__nand3_1 _3141_ (.A(_0221_),
    .B(_0203_),
    .C(_0205_),
    .Y(_0222_));
 sky130_fd_sc_hd__nand2_1 _3142_ (.A(_0220_),
    .B(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__nand2_1 _3143_ (.A(_1311_),
    .B(_1488_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _3144_ (.A(_0223_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__nand3b_1 _3145_ (.A_N(_0224_),
    .B(_0220_),
    .C(_0222_),
    .Y(_0226_));
 sky130_fd_sc_hd__nand2_1 _3146_ (.A(_0225_),
    .B(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _3147_ (.A(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _3148_ (.A(_0142_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21ai_1 _3149_ (.A1(_0229_),
    .A2(_0114_),
    .B1(_0141_),
    .Y(_0230_));
 sky130_fd_sc_hd__or2_1 _3150_ (.A(_0228_),
    .B(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__nand2_1 _3151_ (.A(_0230_),
    .B(_0228_),
    .Y(_0232_));
 sky130_fd_sc_hd__nand2_1 _3152_ (.A(_0231_),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__inv_2 _3153_ (.A(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__nand2_1 _3154_ (.A(_0202_),
    .B(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand3_1 _3155_ (.A(_0199_),
    .B(_0233_),
    .C(_0201_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _3156_ (.A(_0235_),
    .B(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _3157_ (.A(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _3158_ (.A(_0171_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__nand3_1 _3159_ (.A(_0168_),
    .B(_0237_),
    .C(_0170_),
    .Y(_0240_));
 sky130_fd_sc_hd__nand2_1 _3160_ (.A(\datapath.MultiplierAC.PPG0.Y[8] ),
    .B(_1484_),
    .Y(_0241_));
 sky130_fd_sc_hd__xnor2_1 _3161_ (.A(_0154_),
    .B(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__xor2_1 _3162_ (.A(_0155_),
    .B(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__or3_1 _3163_ (.A(_1237_),
    .B(_1510_),
    .C(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__o21ai_1 _3164_ (.A1(_1237_),
    .A2(_1510_),
    .B1(_0243_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand2_1 _3165_ (.A(_0244_),
    .B(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _3166_ (.A(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__a21oi_1 _3167_ (.A1(_0239_),
    .A2(_0240_),
    .B1(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__nand3_1 _3168_ (.A(_0239_),
    .B(_0240_),
    .C(_0247_),
    .Y(_0249_));
 sky130_fd_sc_hd__or2b_1 _3169_ (.A(_0248_),
    .B_N(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _3170_ (.A(_0167_),
    .B(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _3171_ (.A(_0250_),
    .B(_0167_),
    .Y(_0252_));
 sky130_fd_sc_hd__a21oi_1 _3172_ (.A1(_2181_),
    .A2(_2118_),
    .B1(_2180_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand2_1 _3173_ (.A(_1502_),
    .B(_1474_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _3174_ (.A(_1500_),
    .B(_1481_),
    .Y(_0255_));
 sky130_fd_sc_hd__nand2_1 _3175_ (.A(_1498_),
    .B(_1484_),
    .Y(_0256_));
 sky130_fd_sc_hd__nand2_1 _3176_ (.A(_0255_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__o21ai_1 _3177_ (.A1(_1572_),
    .A2(_2126_),
    .B1(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__or2_1 _3178_ (.A(_2128_),
    .B(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_1 _3179_ (.A(_0258_),
    .B(_2128_),
    .Y(_0260_));
 sky130_fd_sc_hd__nand2_1 _3180_ (.A(_0259_),
    .B(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__or2_1 _3181_ (.A(_0254_),
    .B(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__nand2_1 _3182_ (.A(_0261_),
    .B(_0254_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand2_1 _3183_ (.A(_0262_),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__inv_2 _3184_ (.A(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand2_1 _3185_ (.A(_2177_),
    .B(_2174_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_1 _3186_ (.A(_2156_),
    .B(_2153_),
    .Y(_0267_));
 sky130_fd_sc_hd__nand2_1 _3187_ (.A(_2147_),
    .B(_2144_),
    .Y(_0268_));
 sky130_fd_sc_hd__nor2_1 _3188_ (.A(_0255_),
    .B(_0254_),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _3189_ (.A(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__nand2_1 _3190_ (.A(_0255_),
    .B(_0254_),
    .Y(_0271_));
 sky130_fd_sc_hd__nand2_1 _3191_ (.A(_0270_),
    .B(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_2 _3192_ (.A(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand2_1 _3193_ (.A(_2140_),
    .B(_2128_),
    .Y(_0274_));
 sky130_fd_sc_hd__or2_1 _3194_ (.A(_0273_),
    .B(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__nand2_1 _3195_ (.A(_0274_),
    .B(_0273_),
    .Y(_0276_));
 sky130_fd_sc_hd__nand2_1 _3196_ (.A(_0275_),
    .B(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _3197_ (.A(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_2 _3198_ (.A(_0256_),
    .Y(_0279_));
 sky130_fd_sc_hd__nand2_1 _3199_ (.A(_0278_),
    .B(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand2_1 _3200_ (.A(_0277_),
    .B(_0256_),
    .Y(_0281_));
 sky130_fd_sc_hd__nand2_1 _3201_ (.A(_0280_),
    .B(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _3202_ (.A(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2_1 _3203_ (.A(_0268_),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__nand3_1 _3204_ (.A(_2147_),
    .B(_0282_),
    .C(_2144_),
    .Y(_0285_));
 sky130_fd_sc_hd__nand2_1 _3205_ (.A(_0284_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__nand2_1 _3206_ (.A(_1496_),
    .B(_1488_),
    .Y(_0287_));
 sky130_fd_sc_hd__nand2_1 _3207_ (.A(_0286_),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_2 _3208_ (.A(_0287_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand3_1 _3209_ (.A(_0284_),
    .B(_0285_),
    .C(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__nand2_1 _3210_ (.A(_0288_),
    .B(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__inv_2 _3211_ (.A(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__nand2_1 _3212_ (.A(_0267_),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__nand3_1 _3213_ (.A(_2156_),
    .B(_0291_),
    .C(_2153_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand2_1 _3214_ (.A(_0293_),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__nand3_1 _3215_ (.A(_2098_),
    .B(_2099_),
    .C(_2166_),
    .Y(_0296_));
 sky130_fd_sc_hd__o21a_1 _3216_ (.A1(_2094_),
    .A2(_2165_),
    .B1(_2164_),
    .X(_0297_));
 sky130_fd_sc_hd__nand2_1 _3217_ (.A(_0296_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__inv_2 _3218_ (.A(_1492_),
    .Y(_0299_));
 sky130_fd_sc_hd__nor2_1 _3219_ (.A(_1490_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2_1 _3220_ (.A(_0298_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__nand3b_1 _3221_ (.A_N(_0300_),
    .B(_0296_),
    .C(_0297_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2_1 _3222_ (.A(_0301_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__nand2_1 _3223_ (.A(_0303_),
    .B(_0287_),
    .Y(_0304_));
 sky130_fd_sc_hd__nand3_1 _3224_ (.A(_0301_),
    .B(_0302_),
    .C(_0289_),
    .Y(_0305_));
 sky130_fd_sc_hd__nand2_1 _3225_ (.A(_0304_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__a21oi_1 _3226_ (.A1(_2167_),
    .A2(_2168_),
    .B1(_2142_),
    .Y(_0307_));
 sky130_fd_sc_hd__or2_1 _3227_ (.A(_2141_),
    .B(_2169_),
    .X(_0308_));
 sky130_fd_sc_hd__o21ai_1 _3228_ (.A1(_0307_),
    .A2(_2160_),
    .B1(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__xor2_1 _3229_ (.A(_0306_),
    .B(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__nand2_1 _3230_ (.A(_0295_),
    .B(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_2 _3231_ (.A(_0310_),
    .Y(_0312_));
 sky130_fd_sc_hd__nand3_1 _3232_ (.A(_0293_),
    .B(_0312_),
    .C(_0294_),
    .Y(_0313_));
 sky130_fd_sc_hd__nand2_1 _3233_ (.A(_0311_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__inv_2 _3234_ (.A(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand2_1 _3235_ (.A(_0266_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand3_1 _3236_ (.A(_0314_),
    .B(_2177_),
    .C(_2174_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand2_1 _3237_ (.A(_0316_),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _3238_ (.A(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__nor2_1 _3239_ (.A(_0265_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _3240_ (.A(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__nand2_1 _3241_ (.A(_0319_),
    .B(_0265_),
    .Y(_0322_));
 sky130_fd_sc_hd__nand2_1 _3242_ (.A(_0321_),
    .B(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__xor2_1 _3243_ (.A(_0253_),
    .B(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__a32o_1 _3244_ (.A1(_0251_),
    .A2(_1513_),
    .A3(_0252_),
    .B1(_1538_),
    .B2(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__nand2_1 _3245_ (.A(_0325_),
    .B(_1517_),
    .Y(_0326_));
 sky130_fd_sc_hd__nand2_1 _3246_ (.A(_1518_),
    .B(_1500_),
    .Y(_0327_));
 sky130_fd_sc_hd__a21oi_1 _3247_ (.A1(_0326_),
    .A2(_0327_),
    .B1(_1545_),
    .Y(_0026_));
 sky130_fd_sc_hd__nand2_1 _3248_ (.A(_0239_),
    .B(_0235_),
    .Y(_0328_));
 sky130_fd_sc_hd__a22o_1 _3249_ (.A1(_1463_),
    .A2(_1502_),
    .B1(_1466_),
    .B2(_1504_),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _3250_ (.A(_1463_),
    .B(_1504_),
    .Y(_0330_));
 sky130_fd_sc_hd__nor2_1 _3251_ (.A(_0179_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_2 _3252_ (.A(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__nand2_1 _3253_ (.A(_0329_),
    .B(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _3254_ (.A(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__nor2_1 _3255_ (.A(_0087_),
    .B(_0180_),
    .Y(_0335_));
 sky130_fd_sc_hd__o21ai_1 _3256_ (.A1(_0182_),
    .A2(_0091_),
    .B1(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__or2_1 _3257_ (.A(_0334_),
    .B(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__nand2_1 _3258_ (.A(_0336_),
    .B(_0334_),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_1 _3259_ (.A(_0337_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand2_1 _3260_ (.A(_1448_),
    .B(_1500_),
    .Y(_0340_));
 sky130_fd_sc_hd__nand2_1 _3261_ (.A(_0339_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__nand3b_1 _3262_ (.A_N(_0340_),
    .B(_0337_),
    .C(_0338_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _3263_ (.A(_0341_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_2 _3264_ (.A(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__nand2_1 _3265_ (.A(_0192_),
    .B(_0186_),
    .Y(_0345_));
 sky130_fd_sc_hd__xor2_1 _3266_ (.A(_0344_),
    .B(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__nand2_1 _3267_ (.A(_1435_),
    .B(_1498_),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _3268_ (.A(_0346_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__or2_1 _3269_ (.A(_0343_),
    .B(_0345_),
    .X(_0349_));
 sky130_fd_sc_hd__inv_2 _3270_ (.A(_0347_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_1 _3271_ (.A(_0345_),
    .B(_0343_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand3_1 _3272_ (.A(_0349_),
    .B(_0350_),
    .C(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _3273_ (.A(_0348_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand3_1 _3274_ (.A(_2191_),
    .B(_0200_),
    .C(_0109_),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_2 _3275_ (.A(_0104_),
    .Y(_0355_));
 sky130_fd_sc_hd__a21boi_1 _3276_ (.A1(_0355_),
    .A2(_0196_),
    .B1_N(_0197_),
    .Y(_0356_));
 sky130_fd_sc_hd__nand2_1 _3277_ (.A(_0354_),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__or2_1 _3278_ (.A(_0353_),
    .B(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__nand2_1 _3279_ (.A(_0357_),
    .B(_0353_),
    .Y(_0359_));
 sky130_fd_sc_hd__nand2_1 _3280_ (.A(_0358_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__nand2_1 _3281_ (.A(_1311_),
    .B(_1490_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2_1 _3282_ (.A(_0220_),
    .B(_0217_),
    .Y(_0362_));
 sky130_fd_sc_hd__nand2_1 _3283_ (.A(_0216_),
    .B(_0210_),
    .Y(_0363_));
 sky130_fd_sc_hd__a22o_1 _3284_ (.A1(_1379_),
    .A2(_1494_),
    .B1(_1411_),
    .B2(_1496_),
    .X(_0364_));
 sky130_fd_sc_hd__nand2_1 _3285_ (.A(_1379_),
    .B(_1496_),
    .Y(_0365_));
 sky130_fd_sc_hd__nor2_1 _3286_ (.A(_0208_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_2 _3287_ (.A(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__nand2_1 _3288_ (.A(_0364_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__inv_2 _3289_ (.A(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__nand2_1 _3290_ (.A(_0363_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__nand3_1 _3291_ (.A(_0216_),
    .B(_0210_),
    .C(_0368_),
    .Y(_0371_));
 sky130_fd_sc_hd__nand2_1 _3292_ (.A(_0370_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _3293_ (.A(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__nand2_1 _3294_ (.A(_1343_),
    .B(_1492_),
    .Y(_0374_));
 sky130_fd_sc_hd__nand2_1 _3295_ (.A(_0373_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__inv_2 _3296_ (.A(_0374_),
    .Y(_0376_));
 sky130_fd_sc_hd__nand2_1 _3297_ (.A(_0372_),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__nand2_1 _3298_ (.A(_0375_),
    .B(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__nand2_1 _3299_ (.A(_0362_),
    .B(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__inv_2 _3300_ (.A(_0378_),
    .Y(_0380_));
 sky130_fd_sc_hd__nand3_1 _3301_ (.A(_0220_),
    .B(_0380_),
    .C(_0217_),
    .Y(_0381_));
 sky130_fd_sc_hd__nand3b_1 _3302_ (.A_N(_0361_),
    .B(_0379_),
    .C(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_1 _3303_ (.A(_0362_),
    .B(_0380_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand3_1 _3304_ (.A(_0220_),
    .B(_0378_),
    .C(_0217_),
    .Y(_0384_));
 sky130_fd_sc_hd__nand3_1 _3305_ (.A(_0383_),
    .B(_0361_),
    .C(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__and2_1 _3306_ (.A(_0382_),
    .B(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__nand2_1 _3307_ (.A(_0232_),
    .B(_0226_),
    .Y(_0387_));
 sky130_fd_sc_hd__or2_1 _3308_ (.A(_0386_),
    .B(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__nand2_1 _3309_ (.A(_0387_),
    .B(_0386_),
    .Y(_0389_));
 sky130_fd_sc_hd__nand2_1 _3310_ (.A(_0388_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__nand2_1 _3311_ (.A(_0360_),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__inv_2 _3312_ (.A(_0390_),
    .Y(_0392_));
 sky130_fd_sc_hd__nand3_1 _3313_ (.A(_0392_),
    .B(_0358_),
    .C(_0359_),
    .Y(_0393_));
 sky130_fd_sc_hd__nand2_1 _3314_ (.A(_0391_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__inv_2 _3315_ (.A(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__nand2_1 _3316_ (.A(_0328_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__nand3_1 _3317_ (.A(_0239_),
    .B(_0394_),
    .C(_0235_),
    .Y(_0397_));
 sky130_fd_sc_hd__nand2_1 _3318_ (.A(_0396_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__nand2_1 _3319_ (.A(\datapath.MultiplierAC.PPG0.Y[10] ),
    .B(_1482_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _3320_ (.A(\datapath.MultiplierAC.PPG0.Y[9] ),
    .B(_1487_),
    .Y(_0400_));
 sky130_fd_sc_hd__nor2_1 _3321_ (.A(_0241_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__inv_2 _3322_ (.A(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__nand2_1 _3323_ (.A(\datapath.MultiplierAC.PPG0.Y[9] ),
    .B(_1484_),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _3324_ (.A(\datapath.MultiplierAC.PPG0.Y[8] ),
    .B(_1487_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand2_1 _3325_ (.A(_0403_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__nand2_1 _3326_ (.A(_0402_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__a21oi_1 _3327_ (.A1(_2047_),
    .A2(_0241_),
    .B1(_0154_),
    .Y(_0407_));
 sky130_fd_sc_hd__inv_2 _3328_ (.A(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__or2_1 _3329_ (.A(_0406_),
    .B(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__nand2_1 _3330_ (.A(_0408_),
    .B(_0406_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _3331_ (.A(_0409_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__or2_1 _3332_ (.A(_0399_),
    .B(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__nand2_1 _3333_ (.A(_0411_),
    .B(_0399_),
    .Y(_0413_));
 sky130_fd_sc_hd__nand2_1 _3334_ (.A(_0412_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__or2_1 _3335_ (.A(_0414_),
    .B(_0244_),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_1 _3336_ (.A(_0244_),
    .B(_0414_),
    .Y(_0416_));
 sky130_fd_sc_hd__nand2_1 _3337_ (.A(_0415_),
    .B(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__or3_1 _3338_ (.A(_1194_),
    .B(_1510_),
    .C(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__o21ai_1 _3339_ (.A1(_1194_),
    .A2(_1510_),
    .B1(_0417_),
    .Y(_0419_));
 sky130_fd_sc_hd__nand2_1 _3340_ (.A(_0418_),
    .B(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2_1 _3341_ (.A(_0398_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__nand3b_1 _3342_ (.A_N(_0420_),
    .B(_0396_),
    .C(_0397_),
    .Y(_0422_));
 sky130_fd_sc_hd__nand2_1 _3343_ (.A(_0421_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_2 _3344_ (.A(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__o21ai_1 _3345_ (.A1(_0248_),
    .A2(_0167_),
    .B1(_0249_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand2_1 _3346_ (.A(_0424_),
    .B(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__or2_1 _3347_ (.A(_0425_),
    .B(_0424_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _3348_ (.A(_0316_),
    .B(_0313_),
    .Y(_0428_));
 sky130_fd_sc_hd__nand2_1 _3349_ (.A(_0293_),
    .B(_0290_),
    .Y(_0429_));
 sky130_fd_sc_hd__nand2_1 _3350_ (.A(_0284_),
    .B(_0280_),
    .Y(_0430_));
 sky130_fd_sc_hd__nand2_1 _3351_ (.A(_0276_),
    .B(_0270_),
    .Y(_0431_));
 sky130_fd_sc_hd__nand2_1 _3352_ (.A(_1502_),
    .B(_1481_),
    .Y(_0432_));
 sky130_fd_sc_hd__nand2_1 _3353_ (.A(_1504_),
    .B(_1474_),
    .Y(_0433_));
 sky130_fd_sc_hd__nor2_1 _3354_ (.A(_0432_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__inv_2 _3355_ (.A(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__nand2_1 _3356_ (.A(_0432_),
    .B(_0433_),
    .Y(_0436_));
 sky130_fd_sc_hd__nand2_1 _3357_ (.A(_0435_),
    .B(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__inv_2 _3358_ (.A(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__nand2_1 _3359_ (.A(_0431_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__nand3_1 _3360_ (.A(_0276_),
    .B(_0270_),
    .C(_0437_),
    .Y(_0440_));
 sky130_fd_sc_hd__nand2_1 _3361_ (.A(_0439_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__nand2_1 _3362_ (.A(_1500_),
    .B(_1484_),
    .Y(_0442_));
 sky130_fd_sc_hd__nand2_1 _3363_ (.A(_0441_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand3b_1 _3364_ (.A_N(_0442_),
    .B(_0439_),
    .C(_0440_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _3365_ (.A(_0443_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__inv_2 _3366_ (.A(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__nand2_1 _3367_ (.A(_0430_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nand3_1 _3368_ (.A(_0284_),
    .B(_0280_),
    .C(_0445_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand2_1 _3369_ (.A(_0447_),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2_1 _3370_ (.A(_1498_),
    .B(_1487_),
    .Y(_0450_));
 sky130_fd_sc_hd__nand2_1 _3371_ (.A(_0449_),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_2 _3372_ (.A(_0450_),
    .Y(_0452_));
 sky130_fd_sc_hd__nand3_2 _3373_ (.A(_0447_),
    .B(_0452_),
    .C(_0448_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_1 _3374_ (.A(_0451_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_2 _3375_ (.A(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_1 _3376_ (.A(_0429_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__nand3_1 _3377_ (.A(_0293_),
    .B(_0454_),
    .C(_0290_),
    .Y(_0457_));
 sky130_fd_sc_hd__nand2_1 _3378_ (.A(_0456_),
    .B(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_2 _3379_ (.A(_1494_),
    .Y(_0459_));
 sky130_fd_sc_hd__inv_2 _3380_ (.A(_1496_),
    .Y(_0460_));
 sky130_fd_sc_hd__nand2_1 _3381_ (.A(_1496_),
    .B(_1492_),
    .Y(_0461_));
 sky130_fd_sc_hd__nand2_1 _3382_ (.A(_0461_),
    .B(_1490_),
    .Y(_0462_));
 sky130_fd_sc_hd__a21o_1 _3383_ (.A1(_0460_),
    .A2(_0299_),
    .B1(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__o211ai_1 _3384_ (.A1(_0459_),
    .A2(_1657_),
    .B1(_0463_),
    .C1(_0301_),
    .Y(_0464_));
 sky130_fd_sc_hd__or3_1 _3385_ (.A(_0459_),
    .B(_1657_),
    .C(_0463_),
    .X(_0465_));
 sky130_fd_sc_hd__nand2_1 _3386_ (.A(_0464_),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__nand2_1 _3387_ (.A(_1496_),
    .B(_1490_),
    .Y(_0467_));
 sky130_fd_sc_hd__nand2_1 _3388_ (.A(_0466_),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_2 _3389_ (.A(_0467_),
    .Y(_0469_));
 sky130_fd_sc_hd__nand3_1 _3390_ (.A(_0464_),
    .B(_0469_),
    .C(_0465_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2_1 _3391_ (.A(_0468_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__inv_2 _3392_ (.A(_0306_),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_1 _3393_ (.A(_0309_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__nand2_1 _3394_ (.A(_0473_),
    .B(_0305_),
    .Y(_0474_));
 sky130_fd_sc_hd__xor2_1 _3395_ (.A(_0471_),
    .B(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__nand2_1 _3396_ (.A(_0458_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_2 _3397_ (.A(_0475_),
    .Y(_0477_));
 sky130_fd_sc_hd__nand3_1 _3398_ (.A(_0456_),
    .B(_0477_),
    .C(_0457_),
    .Y(_0478_));
 sky130_fd_sc_hd__nand2_1 _3399_ (.A(_0476_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__inv_2 _3400_ (.A(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__nand2_2 _3401_ (.A(_0428_),
    .B(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__nand3_1 _3402_ (.A(_0479_),
    .B(_0316_),
    .C(_0313_),
    .Y(_0482_));
 sky130_fd_sc_hd__nand2_1 _3403_ (.A(_0481_),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__a21oi_1 _3404_ (.A1(_2050_),
    .A2(_0256_),
    .B1(_0255_),
    .Y(_0484_));
 sky130_fd_sc_hd__nor2_1 _3405_ (.A(_1576_),
    .B(_2126_),
    .Y(_0485_));
 sky130_fd_sc_hd__inv_2 _3406_ (.A(_0485_),
    .Y(_0486_));
 sky130_fd_sc_hd__nand2_1 _3407_ (.A(_0442_),
    .B(_0450_),
    .Y(_0487_));
 sky130_fd_sc_hd__and2_1 _3408_ (.A(_0486_),
    .B(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__or2_1 _3409_ (.A(_0484_),
    .B(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nand2_1 _3410_ (.A(_0488_),
    .B(_0484_),
    .Y(_0490_));
 sky130_fd_sc_hd__nand2_1 _3411_ (.A(_0489_),
    .B(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__or2_1 _3412_ (.A(_0432_),
    .B(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_1 _3413_ (.A(_0491_),
    .B(_0432_),
    .Y(_0493_));
 sky130_fd_sc_hd__nand2_1 _3414_ (.A(_0492_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__or2_1 _3415_ (.A(_0262_),
    .B(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__nand2_1 _3416_ (.A(_0494_),
    .B(_0262_),
    .Y(_0496_));
 sky130_fd_sc_hd__nand2_1 _3417_ (.A(_0495_),
    .B(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__or2_1 _3418_ (.A(_0433_),
    .B(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__nand2_1 _3419_ (.A(_0497_),
    .B(_0433_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _3420_ (.A(_0498_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__inv_2 _3421_ (.A(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__nand2_1 _3422_ (.A(_0483_),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__nand3_1 _3423_ (.A(_0481_),
    .B(_0482_),
    .C(_0500_),
    .Y(_0503_));
 sky130_fd_sc_hd__nand2_1 _3424_ (.A(_0502_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__o21ai_1 _3425_ (.A1(_0253_),
    .A2(_0320_),
    .B1(_0322_),
    .Y(_0505_));
 sky130_fd_sc_hd__or2_1 _3426_ (.A(_0504_),
    .B(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__nand2_1 _3427_ (.A(_0505_),
    .B(_0504_),
    .Y(_0507_));
 sky130_fd_sc_hd__and3_1 _3428_ (.A(_0506_),
    .B(_1538_),
    .C(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__a31o_1 _3429_ (.A1(_1513_),
    .A2(_0426_),
    .A3(_0427_),
    .B1(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_1 _3430_ (.A(_0509_),
    .B(_1517_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_1 _3431_ (.A(_1518_),
    .B(_1502_),
    .Y(_0511_));
 sky130_fd_sc_hd__a21oi_1 _3432_ (.A1(_0510_),
    .A2(_0511_),
    .B1(_1545_),
    .Y(_0027_));
 sky130_fd_sc_hd__nand2_1 _3433_ (.A(_0426_),
    .B(_0422_),
    .Y(_0512_));
 sky130_fd_sc_hd__nand2_1 _3434_ (.A(_0396_),
    .B(_0393_),
    .Y(_0513_));
 sky130_fd_sc_hd__or2_1 _3435_ (.A(_0343_),
    .B(_0192_),
    .X(_0514_));
 sky130_fd_sc_hd__nand2_1 _3436_ (.A(_1448_),
    .B(_1502_),
    .Y(_0515_));
 sky130_fd_sc_hd__nand2_1 _3437_ (.A(_1466_),
    .B(\datapath.MultiplierAC.PPG0.X[12] ),
    .Y(_0516_));
 sky130_fd_sc_hd__xnor2_1 _3438_ (.A(_0330_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__nand2_1 _3439_ (.A(_0338_),
    .B(_0332_),
    .Y(_0518_));
 sky130_fd_sc_hd__xor2_1 _3440_ (.A(_0517_),
    .B(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__or2_1 _3441_ (.A(_0515_),
    .B(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__nand2_1 _3442_ (.A(_0519_),
    .B(_0515_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _3443_ (.A(_0520_),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _3444_ (.A(_0342_),
    .B(_0186_),
    .Y(_0523_));
 sky130_fd_sc_hd__nand2_1 _3445_ (.A(_0523_),
    .B(_0341_),
    .Y(_0524_));
 sky130_fd_sc_hd__nand3_1 _3446_ (.A(_0514_),
    .B(_0522_),
    .C(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_2 _3447_ (.A(_0522_),
    .Y(_0526_));
 sky130_fd_sc_hd__o21ai_1 _3448_ (.A1(_0343_),
    .A2(_0192_),
    .B1(_0524_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2_1 _3449_ (.A(_0526_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand2_1 _3450_ (.A(_0525_),
    .B(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand2_1 _3451_ (.A(_1435_),
    .B(_1500_),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _3452_ (.A(_0529_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__nand3b_1 _3453_ (.A_N(_0530_),
    .B(_0525_),
    .C(_0528_),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2_1 _3454_ (.A(_0531_),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__nand2_1 _3455_ (.A(_0346_),
    .B(_0350_),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _3456_ (.A(_0359_),
    .B(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__or2_1 _3457_ (.A(_0533_),
    .B(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__nand2_1 _3458_ (.A(_0535_),
    .B(_0533_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_1 _3459_ (.A(_0536_),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand2_1 _3460_ (.A(_0373_),
    .B(_0376_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _3461_ (.A(_0379_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _3462_ (.A(_1411_),
    .B(_1498_),
    .Y(_0541_));
 sky130_fd_sc_hd__nor2_1 _3463_ (.A(_0365_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_1 _3464_ (.A(_0365_),
    .B(_0541_),
    .Y(_0543_));
 sky130_fd_sc_hd__and2b_1 _3465_ (.A_N(_0542_),
    .B(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__nand2_1 _3466_ (.A(_0370_),
    .B(_0367_),
    .Y(_0545_));
 sky130_fd_sc_hd__or2_1 _3467_ (.A(_0544_),
    .B(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__nand2_1 _3468_ (.A(_0545_),
    .B(_0544_),
    .Y(_0547_));
 sky130_fd_sc_hd__nand2_1 _3469_ (.A(_0546_),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__nand2_1 _3470_ (.A(_1343_),
    .B(_1494_),
    .Y(_0549_));
 sky130_fd_sc_hd__nand2_1 _3471_ (.A(_0548_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__nand3b_1 _3472_ (.A_N(_0549_),
    .B(_0546_),
    .C(_0547_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_1 _3473_ (.A(_0550_),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__inv_2 _3474_ (.A(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__nand2_1 _3475_ (.A(_0540_),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__nand3_1 _3476_ (.A(_0379_),
    .B(_0552_),
    .C(_0539_),
    .Y(_0555_));
 sky130_fd_sc_hd__nand2_1 _3477_ (.A(_0554_),
    .B(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _3478_ (.A(_1311_),
    .B(_1492_),
    .Y(_0557_));
 sky130_fd_sc_hd__nand2_1 _3479_ (.A(_0556_),
    .B(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__nand3b_1 _3480_ (.A_N(_0557_),
    .B(_0554_),
    .C(_0555_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _3481_ (.A(_0558_),
    .B(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__inv_2 _3482_ (.A(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_1 _3483_ (.A(_0389_),
    .B(_0382_),
    .Y(_0562_));
 sky130_fd_sc_hd__or2_1 _3484_ (.A(_0561_),
    .B(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__nand2_1 _3485_ (.A(_0562_),
    .B(_0561_),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2_1 _3486_ (.A(_0563_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__inv_2 _3487_ (.A(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__nand2_1 _3488_ (.A(_0538_),
    .B(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand3_1 _3489_ (.A(_0536_),
    .B(_0565_),
    .C(_0537_),
    .Y(_0568_));
 sky130_fd_sc_hd__nand2_1 _3490_ (.A(_0567_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__inv_2 _3491_ (.A(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_2 _3492_ (.A(_0513_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__nand3_1 _3493_ (.A(_0396_),
    .B(_0569_),
    .C(_0393_),
    .Y(_0572_));
 sky130_fd_sc_hd__nand2_1 _3494_ (.A(_0571_),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__nand2_1 _3495_ (.A(\datapath.MultiplierAC.PPG0.Y[12] ),
    .B(_1475_),
    .Y(_0574_));
 sky130_fd_sc_hd__nand2_1 _3496_ (.A(_0415_),
    .B(_0412_),
    .Y(_0575_));
 sky130_fd_sc_hd__inv_2 _3497_ (.A(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__nand2_1 _3498_ (.A(\datapath.MultiplierAC.PPG0.Y[8] ),
    .B(_1490_),
    .Y(_0577_));
 sky130_fd_sc_hd__or2_1 _3499_ (.A(_0400_),
    .B(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__nand2_1 _3500_ (.A(_0400_),
    .B(_0577_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand2_1 _3501_ (.A(_0578_),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__nand2_1 _3502_ (.A(_0409_),
    .B(_0402_),
    .Y(_0581_));
 sky130_fd_sc_hd__xor2_1 _3503_ (.A(_0580_),
    .B(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__or3_1 _3504_ (.A(_1237_),
    .B(_1636_),
    .C(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__o21ai_1 _3505_ (.A1(_1237_),
    .A2(_1636_),
    .B1(_0582_),
    .Y(_0584_));
 sky130_fd_sc_hd__nand2_1 _3506_ (.A(_0583_),
    .B(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__or2_1 _3507_ (.A(_0576_),
    .B(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__nand2_1 _3508_ (.A(_0585_),
    .B(_0576_),
    .Y(_0587_));
 sky130_fd_sc_hd__nand2_1 _3509_ (.A(_0586_),
    .B(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__nand3b_1 _3510_ (.A_N(_0588_),
    .B(\datapath.MultiplierAC.PPG0.Y[11] ),
    .C(_1482_),
    .Y(_0589_));
 sky130_fd_sc_hd__o21ai_1 _3511_ (.A1(_1194_),
    .A2(_1539_),
    .B1(_0588_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _3512_ (.A(_0589_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__or2_1 _3513_ (.A(_0418_),
    .B(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__nand2_1 _3514_ (.A(_0591_),
    .B(_0418_),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _3515_ (.A(_0592_),
    .B(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__or2_1 _3516_ (.A(_0574_),
    .B(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__nand2_1 _3517_ (.A(_0594_),
    .B(_0574_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _3518_ (.A(_0595_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_1 _3519_ (.A(_0573_),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__inv_2 _3520_ (.A(_0597_),
    .Y(_0599_));
 sky130_fd_sc_hd__nand3_1 _3521_ (.A(_0571_),
    .B(_0572_),
    .C(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__nand2_1 _3522_ (.A(_0598_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__inv_2 _3523_ (.A(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_1 _3524_ (.A(_0512_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__or2_1 _3525_ (.A(_0602_),
    .B(_0512_),
    .X(_0604_));
 sky130_fd_sc_hd__or2_1 _3526_ (.A(_0500_),
    .B(_0483_),
    .X(_0605_));
 sky130_fd_sc_hd__nand2_1 _3527_ (.A(_0507_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _3528_ (.A(_0481_),
    .B(_0478_),
    .Y(_0607_));
 sky130_fd_sc_hd__nand2_1 _3529_ (.A(_0456_),
    .B(_0453_),
    .Y(_0608_));
 sky130_fd_sc_hd__nor2_1 _3530_ (.A(_0282_),
    .B(_0445_),
    .Y(_0609_));
 sky130_fd_sc_hd__nand2_1 _3531_ (.A(_0609_),
    .B(_0268_),
    .Y(_0610_));
 sky130_fd_sc_hd__inv_2 _3532_ (.A(_0280_),
    .Y(_0611_));
 sky130_fd_sc_hd__a21boi_1 _3533_ (.A1(_0611_),
    .A2(_0443_),
    .B1_N(_0444_),
    .Y(_0612_));
 sky130_fd_sc_hd__nand2_1 _3534_ (.A(_0610_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__nand2_1 _3535_ (.A(_0439_),
    .B(_0435_),
    .Y(_0614_));
 sky130_fd_sc_hd__nand2_2 _3536_ (.A(\datapath.MultiplierAC.PPG0.X[12] ),
    .B(_1474_),
    .Y(_0615_));
 sky130_fd_sc_hd__nand2_1 _3537_ (.A(_1504_),
    .B(_1482_),
    .Y(_0616_));
 sky130_fd_sc_hd__nor2_1 _3538_ (.A(_0615_),
    .B(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__nand2_1 _3539_ (.A(_0615_),
    .B(_0616_),
    .Y(_0618_));
 sky130_fd_sc_hd__inv_2 _3540_ (.A(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__nor2_1 _3541_ (.A(_0617_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__nand2_1 _3542_ (.A(_0614_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__inv_2 _3543_ (.A(_0620_),
    .Y(_0622_));
 sky130_fd_sc_hd__nand3_1 _3544_ (.A(_0439_),
    .B(_0435_),
    .C(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2_1 _3545_ (.A(_0621_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _3546_ (.A(_1502_),
    .B(_1485_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand2_1 _3547_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__nand3b_2 _3548_ (.A_N(_0625_),
    .B(_0621_),
    .C(_0623_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2_1 _3549_ (.A(_0626_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__inv_2 _3550_ (.A(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__nand2_1 _3551_ (.A(_0613_),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__nand3_1 _3552_ (.A(_0610_),
    .B(_0628_),
    .C(_0612_),
    .Y(_0631_));
 sky130_fd_sc_hd__nand2_1 _3553_ (.A(_0630_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__nand2_1 _3554_ (.A(_1500_),
    .B(_1487_),
    .Y(_0633_));
 sky130_fd_sc_hd__nand2_1 _3555_ (.A(_0632_),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__nand3b_1 _3556_ (.A_N(_0633_),
    .B(_0630_),
    .C(_0631_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand2_1 _3557_ (.A(_0634_),
    .B(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__inv_2 _3558_ (.A(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__nand2_1 _3559_ (.A(_0608_),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__nand3_1 _3560_ (.A(_0456_),
    .B(_0453_),
    .C(_0636_),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_1 _3561_ (.A(_0638_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__nor2_1 _3562_ (.A(_1492_),
    .B(_0469_),
    .Y(_0641_));
 sky130_fd_sc_hd__nand2_1 _3563_ (.A(_0641_),
    .B(_1494_),
    .Y(_0642_));
 sky130_fd_sc_hd__o21ai_1 _3564_ (.A1(_1496_),
    .A2(_1494_),
    .B1(_1709_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand2_1 _3565_ (.A(_1498_),
    .B(\datapath.MultiplierAC.PPG0.X[4] ),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_1 _3566_ (.A(_0461_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__o21ai_1 _3567_ (.A1(_1708_),
    .A2(_2059_),
    .B1(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__or2_1 _3568_ (.A(_0643_),
    .B(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__nand2_1 _3569_ (.A(_0646_),
    .B(_0643_),
    .Y(_0648_));
 sky130_fd_sc_hd__nand2_1 _3570_ (.A(_0647_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__xnor2_1 _3571_ (.A(_0642_),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__or2_1 _3572_ (.A(_0461_),
    .B(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__nand2_1 _3573_ (.A(_0650_),
    .B(_0461_),
    .Y(_0652_));
 sky130_fd_sc_hd__nand2_1 _3574_ (.A(_0651_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__inv_2 _3575_ (.A(_0471_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand2_1 _3576_ (.A(_0474_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__nand2_1 _3577_ (.A(_0655_),
    .B(_0470_),
    .Y(_0656_));
 sky130_fd_sc_hd__xor2_1 _3578_ (.A(_0653_),
    .B(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__nand2_1 _3579_ (.A(_0640_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__inv_2 _3580_ (.A(_0657_),
    .Y(_0659_));
 sky130_fd_sc_hd__nand3_2 _3581_ (.A(_0638_),
    .B(_0659_),
    .C(_0639_),
    .Y(_0660_));
 sky130_fd_sc_hd__nand2_1 _3582_ (.A(_0658_),
    .B(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__inv_2 _3583_ (.A(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__nand2_1 _3584_ (.A(_0607_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__nand3_1 _3585_ (.A(_0661_),
    .B(_0481_),
    .C(_0478_),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _3586_ (.A(_0663_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__nor2_1 _3587_ (.A(_0633_),
    .B(_0644_),
    .Y(_0666_));
 sky130_fd_sc_hd__inv_2 _3588_ (.A(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__nand2_1 _3589_ (.A(_0633_),
    .B(_0644_),
    .Y(_0668_));
 sky130_fd_sc_hd__and2_1 _3590_ (.A(_0667_),
    .B(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__nand2_1 _3591_ (.A(_0490_),
    .B(_0486_),
    .Y(_0670_));
 sky130_fd_sc_hd__or2_1 _3592_ (.A(_0669_),
    .B(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__nand2_1 _3593_ (.A(_0670_),
    .B(_0669_),
    .Y(_0672_));
 sky130_fd_sc_hd__nand2_1 _3594_ (.A(_0671_),
    .B(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__or2_1 _3595_ (.A(_0625_),
    .B(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__nand2_1 _3596_ (.A(_0673_),
    .B(_0625_),
    .Y(_0675_));
 sky130_fd_sc_hd__nand2_1 _3597_ (.A(_0674_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__inv_2 _3598_ (.A(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand2_1 _3599_ (.A(_0495_),
    .B(_0492_),
    .Y(_0678_));
 sky130_fd_sc_hd__or2_1 _3600_ (.A(_0677_),
    .B(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__nand2_1 _3601_ (.A(_0678_),
    .B(_0677_),
    .Y(_0680_));
 sky130_fd_sc_hd__nand2_1 _3602_ (.A(_0679_),
    .B(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__or2_1 _3603_ (.A(_0616_),
    .B(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__nand2_1 _3604_ (.A(_0681_),
    .B(_0616_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _3605_ (.A(_0682_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__or2_1 _3606_ (.A(_0498_),
    .B(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__nand2_1 _3607_ (.A(_0684_),
    .B(_0498_),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_1 _3608_ (.A(_0685_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__inv_2 _3609_ (.A(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__inv_2 _3610_ (.A(_0615_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2_1 _3611_ (.A(_0688_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__nand2_1 _3612_ (.A(_0687_),
    .B(_0615_),
    .Y(_0691_));
 sky130_fd_sc_hd__nand2_1 _3613_ (.A(_0690_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_1 _3614_ (.A(_0665_),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__nand3b_1 _3615_ (.A_N(_0692_),
    .B(_0663_),
    .C(_0664_),
    .Y(_0694_));
 sky130_fd_sc_hd__nand2_1 _3616_ (.A(_0693_),
    .B(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__inv_2 _3617_ (.A(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__or2_1 _3618_ (.A(_0606_),
    .B(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__nand2_1 _3619_ (.A(_0696_),
    .B(_0606_),
    .Y(_0698_));
 sky130_fd_sc_hd__and3_1 _3620_ (.A(_0697_),
    .B(_1538_),
    .C(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__a31o_1 _3621_ (.A1(_1513_),
    .A2(_0603_),
    .A3(_0604_),
    .B1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__nand2_1 _3622_ (.A(_0700_),
    .B(_1517_),
    .Y(_0701_));
 sky130_fd_sc_hd__nand2_1 _3623_ (.A(_1518_),
    .B(_1504_),
    .Y(_0702_));
 sky130_fd_sc_hd__a21oi_1 _3624_ (.A1(_0701_),
    .A2(_0702_),
    .B1(_1545_),
    .Y(_0028_));
 sky130_fd_sc_hd__nand2_1 _3625_ (.A(_0663_),
    .B(_0660_),
    .Y(_0703_));
 sky130_fd_sc_hd__nor2_1 _3626_ (.A(_0454_),
    .B(_0636_),
    .Y(_0704_));
 sky130_fd_sc_hd__nand2_1 _3627_ (.A(_0704_),
    .B(_0429_),
    .Y(_0705_));
 sky130_fd_sc_hd__inv_2 _3628_ (.A(_0453_),
    .Y(_0706_));
 sky130_fd_sc_hd__a21boi_1 _3629_ (.A1(_0634_),
    .A2(_0706_),
    .B1_N(_0635_),
    .Y(_0707_));
 sky130_fd_sc_hd__nand2_1 _3630_ (.A(_0705_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__nand2_1 _3631_ (.A(_0630_),
    .B(_0627_),
    .Y(_0709_));
 sky130_fd_sc_hd__a22o_1 _3632_ (.A1(\datapath.MultiplierAC.PPG0.X[13] ),
    .A2(_1475_),
    .B1(\datapath.MultiplierAC.PPG0.X[12] ),
    .B2(_1482_),
    .X(_0710_));
 sky130_fd_sc_hd__nand2_1 _3633_ (.A(\datapath.MultiplierAC.PPG0.X[13] ),
    .B(_1482_),
    .Y(_0711_));
 sky130_fd_sc_hd__nor2_1 _3634_ (.A(_0615_),
    .B(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__inv_2 _3635_ (.A(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__nand2_1 _3636_ (.A(_0710_),
    .B(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__inv_2 _3637_ (.A(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__and4_1 _3638_ (.A(_2133_),
    .B(_0273_),
    .C(_0438_),
    .D(_0620_),
    .X(_0716_));
 sky130_fd_sc_hd__nand2_1 _3639_ (.A(_0716_),
    .B(_2138_),
    .Y(_0717_));
 sky130_fd_sc_hd__a21oi_1 _3640_ (.A1(_2050_),
    .A2(_0254_),
    .B1(_0255_),
    .Y(_0718_));
 sky130_fd_sc_hd__a311o_1 _3641_ (.A1(_0718_),
    .A2(_0436_),
    .A3(_0618_),
    .B1(_0434_),
    .C1(_0617_),
    .X(_0719_));
 sky130_fd_sc_hd__inv_2 _3642_ (.A(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__nand2_1 _3643_ (.A(_0717_),
    .B(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__or2_1 _3644_ (.A(_0715_),
    .B(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__nand2_1 _3645_ (.A(_0721_),
    .B(_0715_),
    .Y(_0723_));
 sky130_fd_sc_hd__nand2_1 _3646_ (.A(_0722_),
    .B(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__nand2_1 _3647_ (.A(_1504_),
    .B(_1485_),
    .Y(_0725_));
 sky130_fd_sc_hd__nand2_1 _3648_ (.A(_0724_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand3b_1 _3649_ (.A_N(_0725_),
    .B(_0722_),
    .C(_0723_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_1 _3650_ (.A(_0726_),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__inv_2 _3651_ (.A(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__nand2_1 _3652_ (.A(_0709_),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__nand3_1 _3653_ (.A(_0630_),
    .B(_0627_),
    .C(_0728_),
    .Y(_0731_));
 sky130_fd_sc_hd__nand2_1 _3654_ (.A(_0730_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__nand2_1 _3655_ (.A(_1502_),
    .B(_1488_),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_1 _3656_ (.A(_0732_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand3b_1 _3657_ (.A_N(_0733_),
    .B(_0730_),
    .C(_0731_),
    .Y(_0735_));
 sky130_fd_sc_hd__nand2_1 _3658_ (.A(_0734_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__inv_2 _3659_ (.A(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _3660_ (.A(_0708_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__nand3_1 _3661_ (.A(_0705_),
    .B(_0736_),
    .C(_0707_),
    .Y(_0739_));
 sky130_fd_sc_hd__nand2_1 _3662_ (.A(_0738_),
    .B(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__inv_2 _3663_ (.A(_0653_),
    .Y(_0741_));
 sky130_fd_sc_hd__nand2_1 _3664_ (.A(_0656_),
    .B(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__nand2_1 _3665_ (.A(_0742_),
    .B(_0651_),
    .Y(_0743_));
 sky130_fd_sc_hd__a21o_1 _3666_ (.A1(_0649_),
    .A2(_0641_),
    .B1(_0459_),
    .X(_0744_));
 sky130_fd_sc_hd__a22o_1 _3667_ (.A1(_1500_),
    .A2(_1490_),
    .B1(_1498_),
    .B2(_1492_),
    .X(_0745_));
 sky130_fd_sc_hd__nand2_1 _3668_ (.A(_1500_),
    .B(\datapath.MultiplierAC.PPG0.X[5] ),
    .Y(_0746_));
 sky130_fd_sc_hd__or2_1 _3669_ (.A(_0644_),
    .B(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__nand2_1 _3670_ (.A(_0745_),
    .B(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__o21a_1 _3671_ (.A1(_1708_),
    .A2(_2059_),
    .B1(_0647_),
    .X(_0749_));
 sky130_fd_sc_hd__or2_1 _3672_ (.A(_0748_),
    .B(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__nand2_1 _3673_ (.A(_0749_),
    .B(_0748_),
    .Y(_0751_));
 sky130_fd_sc_hd__nand2_1 _3674_ (.A(_0750_),
    .B(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__or2_1 _3675_ (.A(_1929_),
    .B(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__nand2_1 _3676_ (.A(_0752_),
    .B(_1929_),
    .Y(_0754_));
 sky130_fd_sc_hd__nand2_1 _3677_ (.A(_0753_),
    .B(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__or2_1 _3678_ (.A(_0744_),
    .B(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__nand2_1 _3679_ (.A(_0755_),
    .B(_0744_),
    .Y(_0757_));
 sky130_fd_sc_hd__nand2_1 _3680_ (.A(_0756_),
    .B(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__nor2_1 _3681_ (.A(_1929_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__inv_2 _3682_ (.A(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _3683_ (.A(_0758_),
    .B(_1929_),
    .Y(_0761_));
 sky130_fd_sc_hd__nand2_1 _3684_ (.A(_0760_),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__inv_2 _3685_ (.A(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__nand2_1 _3686_ (.A(_0743_),
    .B(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__nand3_1 _3687_ (.A(_0742_),
    .B(_0651_),
    .C(_0762_),
    .Y(_0765_));
 sky130_fd_sc_hd__nand2_1 _3688_ (.A(_0764_),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__nand2_1 _3689_ (.A(_0740_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__inv_2 _3690_ (.A(_0766_),
    .Y(_0768_));
 sky130_fd_sc_hd__nand3_1 _3691_ (.A(_0768_),
    .B(_0738_),
    .C(_0739_),
    .Y(_0769_));
 sky130_fd_sc_hd__nand2_1 _3692_ (.A(_0767_),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__inv_2 _3693_ (.A(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__nand2_1 _3694_ (.A(_0703_),
    .B(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__nand3_1 _3695_ (.A(_0663_),
    .B(_0660_),
    .C(_0770_),
    .Y(_0773_));
 sky130_fd_sc_hd__nand2_1 _3696_ (.A(_0772_),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__nand2_1 _3697_ (.A(_0680_),
    .B(_0674_),
    .Y(_0775_));
 sky130_fd_sc_hd__nand2_1 _3698_ (.A(_0672_),
    .B(_0667_),
    .Y(_0776_));
 sky130_fd_sc_hd__inv_2 _3699_ (.A(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__or2_1 _3700_ (.A(_0748_),
    .B(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__nand2_1 _3701_ (.A(_0777_),
    .B(_0748_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2_1 _3702_ (.A(_0778_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__or2_1 _3703_ (.A(_0733_),
    .B(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__nand2_1 _3704_ (.A(_0780_),
    .B(_0733_),
    .Y(_0782_));
 sky130_fd_sc_hd__nand2_1 _3705_ (.A(_0781_),
    .B(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__inv_2 _3706_ (.A(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__or2_1 _3707_ (.A(_0775_),
    .B(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__nand2_1 _3708_ (.A(_0784_),
    .B(_0775_),
    .Y(_0786_));
 sky130_fd_sc_hd__nand2_1 _3709_ (.A(_0785_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__or2_1 _3710_ (.A(_0725_),
    .B(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_1 _3711_ (.A(_0787_),
    .B(_0725_),
    .Y(_0789_));
 sky130_fd_sc_hd__nand2_1 _3712_ (.A(_0788_),
    .B(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__inv_2 _3713_ (.A(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand2_1 _3714_ (.A(_0685_),
    .B(_0682_),
    .Y(_0792_));
 sky130_fd_sc_hd__or2_1 _3715_ (.A(_0791_),
    .B(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__nand2_1 _3716_ (.A(_0792_),
    .B(_0791_),
    .Y(_0794_));
 sky130_fd_sc_hd__a21o_1 _3717_ (.A1(_0793_),
    .A2(_0794_),
    .B1(_0715_),
    .X(_0795_));
 sky130_fd_sc_hd__nand3_1 _3718_ (.A(_0793_),
    .B(_0715_),
    .C(_0794_),
    .Y(_0796_));
 sky130_fd_sc_hd__nand2_1 _3719_ (.A(_0795_),
    .B(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__inv_2 _3720_ (.A(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__inv_2 _3721_ (.A(_0690_),
    .Y(_0799_));
 sky130_fd_sc_hd__nand2_1 _3722_ (.A(_0798_),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand2_1 _3723_ (.A(_0797_),
    .B(_0690_),
    .Y(_0801_));
 sky130_fd_sc_hd__nand2_1 _3724_ (.A(_0800_),
    .B(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__nand2_1 _3725_ (.A(_0774_),
    .B(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__inv_2 _3726_ (.A(_0802_),
    .Y(_0804_));
 sky130_fd_sc_hd__nand3_1 _3727_ (.A(_0772_),
    .B(_0773_),
    .C(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__nand2_1 _3728_ (.A(_0803_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__nand2_1 _3729_ (.A(_0698_),
    .B(_0694_),
    .Y(_0807_));
 sky130_fd_sc_hd__inv_2 _3730_ (.A(_0806_),
    .Y(_0808_));
 sky130_fd_sc_hd__nand2_1 _3731_ (.A(_0807_),
    .B(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__nand2_1 _3732_ (.A(_0809_),
    .B(_1538_),
    .Y(_0810_));
 sky130_fd_sc_hd__a31o_1 _3733_ (.A1(_0694_),
    .A2(_0698_),
    .A3(_0806_),
    .B1(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__nand2_1 _3734_ (.A(\datapath.MultiplierAC.PPG0.Y[10] ),
    .B(_1488_),
    .Y(_0812_));
 sky130_fd_sc_hd__a22o_1 _3735_ (.A1(\datapath.MultiplierAC.PPG0.Y[9] ),
    .A2(_1490_),
    .B1(\datapath.MultiplierAC.PPG0.Y[8] ),
    .B2(_1492_),
    .X(_0813_));
 sky130_fd_sc_hd__nand2_1 _3736_ (.A(\datapath.MultiplierAC.PPG0.Y[9] ),
    .B(_1492_),
    .Y(_0814_));
 sky130_fd_sc_hd__nor2_1 _3737_ (.A(_0577_),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__inv_2 _3738_ (.A(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__nand2_1 _3739_ (.A(_0813_),
    .B(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__and2_1 _3740_ (.A(_0578_),
    .B(_0402_),
    .X(_0818_));
 sky130_fd_sc_hd__inv_2 _3741_ (.A(_0579_),
    .Y(_0819_));
 sky130_fd_sc_hd__a21oi_1 _3742_ (.A1(_0409_),
    .A2(_0818_),
    .B1(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__inv_2 _3743_ (.A(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__or2_1 _3744_ (.A(_0817_),
    .B(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__nand2_1 _3745_ (.A(_0821_),
    .B(_0817_),
    .Y(_0823_));
 sky130_fd_sc_hd__nand2_1 _3746_ (.A(_0822_),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__or2_1 _3747_ (.A(_0812_),
    .B(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__nand2_1 _3748_ (.A(_0824_),
    .B(_0812_),
    .Y(_0826_));
 sky130_fd_sc_hd__and2_1 _3749_ (.A(_0825_),
    .B(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__nand2_1 _3750_ (.A(_0586_),
    .B(_0583_),
    .Y(_0828_));
 sky130_fd_sc_hd__or2_1 _3751_ (.A(_0827_),
    .B(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__nand2_1 _3752_ (.A(_0828_),
    .B(_0827_),
    .Y(_0830_));
 sky130_fd_sc_hd__nand2_1 _3753_ (.A(_0829_),
    .B(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__or3_1 _3754_ (.A(_1194_),
    .B(_1636_),
    .C(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__o21ai_1 _3755_ (.A1(_1194_),
    .A2(_1636_),
    .B1(_0831_),
    .Y(_0833_));
 sky130_fd_sc_hd__nand2_1 _3756_ (.A(_0592_),
    .B(_0589_),
    .Y(_0834_));
 sky130_fd_sc_hd__a21o_1 _3757_ (.A1(_0832_),
    .A2(_0833_),
    .B1(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__nand3_1 _3758_ (.A(_0832_),
    .B(_0834_),
    .C(_0833_),
    .Y(_0836_));
 sky130_fd_sc_hd__nand2_1 _3759_ (.A(_0835_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__inv_2 _3760_ (.A(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__a22o_1 _3761_ (.A1(\datapath.MultiplierAC.PPG0.Y[13] ),
    .A2(_1475_),
    .B1(\datapath.MultiplierAC.PPG0.Y[12] ),
    .B2(_1482_),
    .X(_0839_));
 sky130_fd_sc_hd__nand2_1 _3762_ (.A(\datapath.MultiplierAC.PPG0.Y[13] ),
    .B(_1482_),
    .Y(_0840_));
 sky130_fd_sc_hd__nor2_1 _3763_ (.A(_0574_),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__inv_2 _3764_ (.A(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__nand2_1 _3765_ (.A(_0839_),
    .B(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__inv_2 _3766_ (.A(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__nand2_1 _3767_ (.A(_0838_),
    .B(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__nand2_1 _3768_ (.A(_0837_),
    .B(_0843_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _3769_ (.A(_0845_),
    .B(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__nand2_1 _3770_ (.A(_0847_),
    .B(_0595_),
    .Y(_0848_));
 sky130_fd_sc_hd__inv_2 _3771_ (.A(_0595_),
    .Y(_0849_));
 sky130_fd_sc_hd__nand3_1 _3772_ (.A(_0845_),
    .B(_0846_),
    .C(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _3773_ (.A(_0848_),
    .B(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__nand2_1 _3774_ (.A(_0571_),
    .B(_0567_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand2_1 _3775_ (.A(_0532_),
    .B(_0534_),
    .Y(_0853_));
 sky130_fd_sc_hd__nand2_1 _3776_ (.A(_0853_),
    .B(_0531_),
    .Y(_0854_));
 sky130_fd_sc_hd__o21ai_1 _3777_ (.A1(_0533_),
    .A2(_0359_),
    .B1(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__a22o_1 _3778_ (.A1(_1463_),
    .A2(\datapath.MultiplierAC.PPG0.X[12] ),
    .B1(_1466_),
    .B2(\datapath.MultiplierAC.PPG0.X[13] ),
    .X(_0856_));
 sky130_fd_sc_hd__nand2_1 _3779_ (.A(_1463_),
    .B(\datapath.MultiplierAC.PPG0.X[13] ),
    .Y(_0857_));
 sky130_fd_sc_hd__or2_1 _3780_ (.A(_0516_),
    .B(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__and2_1 _3781_ (.A(_0856_),
    .B(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__nor2_1 _3782_ (.A(_0517_),
    .B(_0333_),
    .Y(_0860_));
 sky130_fd_sc_hd__nand2_1 _3783_ (.A(_0336_),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__a21o_1 _3784_ (.A1(_0179_),
    .A2(_0516_),
    .B1(_0330_),
    .X(_0862_));
 sky130_fd_sc_hd__nand2_1 _3785_ (.A(_0861_),
    .B(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__or2_1 _3786_ (.A(_0859_),
    .B(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__nand2_1 _3787_ (.A(_0863_),
    .B(_0859_),
    .Y(_0865_));
 sky130_fd_sc_hd__nand2_1 _3788_ (.A(_0864_),
    .B(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__nand2_1 _3789_ (.A(_1448_),
    .B(_1504_),
    .Y(_0867_));
 sky130_fd_sc_hd__nand2_1 _3790_ (.A(_0866_),
    .B(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__nand3b_1 _3791_ (.A_N(_0867_),
    .B(_0864_),
    .C(_0865_),
    .Y(_0869_));
 sky130_fd_sc_hd__nand2_1 _3792_ (.A(_0868_),
    .B(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__nand2_1 _3793_ (.A(_0528_),
    .B(_0520_),
    .Y(_0871_));
 sky130_fd_sc_hd__xnor2_1 _3794_ (.A(_0870_),
    .B(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__nand2_1 _3795_ (.A(_1435_),
    .B(_1502_),
    .Y(_0873_));
 sky130_fd_sc_hd__inv_2 _3796_ (.A(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__nand2_1 _3797_ (.A(_0872_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__or2_1 _3798_ (.A(_0870_),
    .B(_0871_),
    .X(_0876_));
 sky130_fd_sc_hd__nand2_1 _3799_ (.A(_0871_),
    .B(_0870_),
    .Y(_0877_));
 sky130_fd_sc_hd__nand3_1 _3800_ (.A(_0876_),
    .B(_0873_),
    .C(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__nand2_1 _3801_ (.A(_0875_),
    .B(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__nand2b_1 _3802_ (.A_N(_0855_),
    .B(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2b_1 _3803_ (.A_N(_0879_),
    .B(_0855_),
    .Y(_0881_));
 sky130_fd_sc_hd__nand2_1 _3804_ (.A(_0880_),
    .B(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__nand2_1 _3805_ (.A(_0564_),
    .B(_0559_),
    .Y(_0883_));
 sky130_fd_sc_hd__nand2_1 _3806_ (.A(_1311_),
    .B(_1494_),
    .Y(_0884_));
 sky130_fd_sc_hd__nand2_1 _3807_ (.A(_0554_),
    .B(_0551_),
    .Y(_0885_));
 sky130_fd_sc_hd__inv_2 _3808_ (.A(_1500_),
    .Y(_0886_));
 sky130_fd_sc_hd__or3_1 _3809_ (.A(_1387_),
    .B(_0886_),
    .C(_0541_),
    .X(_0887_));
 sky130_fd_sc_hd__a22o_1 _3810_ (.A1(_1379_),
    .A2(_1498_),
    .B1(_1411_),
    .B2(_1500_),
    .X(_0888_));
 sky130_fd_sc_hd__and2_1 _3811_ (.A(_0887_),
    .B(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__and4_1 _3812_ (.A(_0126_),
    .B(_0369_),
    .C(_0213_),
    .D(_0544_),
    .X(_0890_));
 sky130_fd_sc_hd__a21oi_1 _3813_ (.A1(_2016_),
    .A2(_0208_),
    .B1(_0121_),
    .Y(_0891_));
 sky130_fd_sc_hd__a311o_1 _3814_ (.A1(_0364_),
    .A2(_0891_),
    .A3(_0543_),
    .B1(_0366_),
    .C1(_0542_),
    .X(_0892_));
 sky130_fd_sc_hd__a21o_1 _3815_ (.A1(_0119_),
    .A2(_0890_),
    .B1(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__or2_1 _3816_ (.A(_0889_),
    .B(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__nand2_1 _3817_ (.A(_0893_),
    .B(_0889_),
    .Y(_0895_));
 sky130_fd_sc_hd__nand2_1 _3818_ (.A(_0894_),
    .B(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__inv_2 _3819_ (.A(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__nand2_1 _3820_ (.A(_1343_),
    .B(_1496_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_1 _3821_ (.A(_0897_),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__inv_2 _3822_ (.A(_0898_),
    .Y(_0900_));
 sky130_fd_sc_hd__nand2_1 _3823_ (.A(_0896_),
    .B(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__nand2_1 _3824_ (.A(_0899_),
    .B(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__nand2_1 _3825_ (.A(_0885_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__inv_2 _3826_ (.A(_0902_),
    .Y(_0904_));
 sky130_fd_sc_hd__nand3_1 _3827_ (.A(_0554_),
    .B(_0551_),
    .C(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__nand3b_1 _3828_ (.A_N(_0884_),
    .B(_0903_),
    .C(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__nand2_1 _3829_ (.A(_0885_),
    .B(_0904_),
    .Y(_0907_));
 sky130_fd_sc_hd__nand3_1 _3830_ (.A(_0554_),
    .B(_0551_),
    .C(_0902_),
    .Y(_0908_));
 sky130_fd_sc_hd__nand3_1 _3831_ (.A(_0907_),
    .B(_0908_),
    .C(_0884_),
    .Y(_0909_));
 sky130_fd_sc_hd__nand2_1 _3832_ (.A(_0906_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__inv_2 _3833_ (.A(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__nand2_1 _3834_ (.A(_0883_),
    .B(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__nand3_1 _3835_ (.A(_0910_),
    .B(_0564_),
    .C(_0559_),
    .Y(_0913_));
 sky130_fd_sc_hd__nand2_1 _3836_ (.A(_0912_),
    .B(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__nand2_1 _3837_ (.A(_0882_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__nand3b_1 _3838_ (.A_N(_0914_),
    .B(_0880_),
    .C(_0881_),
    .Y(_0916_));
 sky130_fd_sc_hd__nand2_1 _3839_ (.A(_0915_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__inv_2 _3840_ (.A(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__nand2_1 _3841_ (.A(_0852_),
    .B(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__nand3_1 _3842_ (.A(_0571_),
    .B(_0567_),
    .C(_0917_),
    .Y(_0920_));
 sky130_fd_sc_hd__nand3b_1 _3843_ (.A_N(_0851_),
    .B(_0919_),
    .C(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__nand2_1 _3844_ (.A(_0852_),
    .B(_0917_),
    .Y(_0922_));
 sky130_fd_sc_hd__nand3_1 _3845_ (.A(_0571_),
    .B(_0918_),
    .C(_0567_),
    .Y(_0923_));
 sky130_fd_sc_hd__nand3_1 _3846_ (.A(_0922_),
    .B(_0923_),
    .C(_0851_),
    .Y(_0924_));
 sky130_fd_sc_hd__nand2_1 _3847_ (.A(_0921_),
    .B(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__inv_2 _3848_ (.A(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__nand2_1 _3849_ (.A(_0603_),
    .B(_0600_),
    .Y(_0927_));
 sky130_fd_sc_hd__or2_1 _3850_ (.A(_0926_),
    .B(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__nand2_1 _3851_ (.A(_0927_),
    .B(_0926_),
    .Y(_0929_));
 sky130_fd_sc_hd__nand3_1 _3852_ (.A(_0928_),
    .B(_1513_),
    .C(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__o21ai_1 _3853_ (.A1(_1517_),
    .A2(\datapath.MultiplierAC.PPG0.X[12] ),
    .B1(_1067_),
    .Y(_0931_));
 sky130_fd_sc_hd__a31oi_1 _3854_ (.A1(_0811_),
    .A2(_0930_),
    .A3(_1517_),
    .B1(_0931_),
    .Y(_0029_));
 sky130_fd_sc_hd__nand2_1 _3855_ (.A(_0929_),
    .B(_0921_),
    .Y(_0932_));
 sky130_fd_sc_hd__or2_1 _3856_ (.A(_0917_),
    .B(_0571_),
    .X(_0933_));
 sky130_fd_sc_hd__nand2_1 _3857_ (.A(_0881_),
    .B(_0875_),
    .Y(_0934_));
 sky130_fd_sc_hd__inv_2 _3858_ (.A(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__inv_2 _3859_ (.A(\datapath.MultiplierAC.PPG0.X[12] ),
    .Y(_0936_));
 sky130_fd_sc_hd__nand2_1 _3860_ (.A(_1466_),
    .B(\datapath.MultiplierAC.PPG0.X[14] ),
    .Y(_0937_));
 sky130_fd_sc_hd__xnor2_1 _3861_ (.A(_0857_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__nand2_1 _3862_ (.A(_0865_),
    .B(_0858_),
    .Y(_0939_));
 sky130_fd_sc_hd__xor2_1 _3863_ (.A(_0938_),
    .B(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__or3_1 _3864_ (.A(_1457_),
    .B(_0936_),
    .C(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__o21ai_1 _3865_ (.A1(_1457_),
    .A2(_0936_),
    .B1(_0940_),
    .Y(_0942_));
 sky130_fd_sc_hd__nor2_1 _3866_ (.A(_0870_),
    .B(_0522_),
    .Y(_0943_));
 sky130_fd_sc_hd__o21ai_1 _3867_ (.A1(_0520_),
    .A2(_0870_),
    .B1(_0869_),
    .Y(_0944_));
 sky130_fd_sc_hd__a21o_1 _3868_ (.A1(_0943_),
    .A2(_0527_),
    .B1(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__a21o_1 _3869_ (.A1(_0941_),
    .A2(_0942_),
    .B1(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__nand3_1 _3870_ (.A(_0945_),
    .B(_0941_),
    .C(_0942_),
    .Y(_0947_));
 sky130_fd_sc_hd__nand2_1 _3871_ (.A(_0946_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__nand2_1 _3872_ (.A(_1435_),
    .B(_1504_),
    .Y(_0949_));
 sky130_fd_sc_hd__nand2_1 _3873_ (.A(_0948_),
    .B(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__nand3b_1 _3874_ (.A_N(_0949_),
    .B(_0946_),
    .C(_0947_),
    .Y(_0951_));
 sky130_fd_sc_hd__nand2_1 _3875_ (.A(_0950_),
    .B(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__inv_2 _3876_ (.A(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__nand2_1 _3877_ (.A(_0935_),
    .B(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__nand2_1 _3878_ (.A(_0934_),
    .B(_0952_),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2_1 _3879_ (.A(_0954_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__nand2_1 _3880_ (.A(_0897_),
    .B(_0900_),
    .Y(_0957_));
 sky130_fd_sc_hd__nand2_1 _3881_ (.A(_0903_),
    .B(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__nand2_1 _3882_ (.A(_1411_),
    .B(_1502_),
    .Y(_0959_));
 sky130_fd_sc_hd__nor3_1 _3883_ (.A(_1387_),
    .B(_0886_),
    .C(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__inv_2 _3884_ (.A(_0960_),
    .Y(_0961_));
 sky130_fd_sc_hd__o21ai_1 _3885_ (.A1(_1387_),
    .A2(_0886_),
    .B1(_0959_),
    .Y(_0962_));
 sky130_fd_sc_hd__nand2_1 _3886_ (.A(_0961_),
    .B(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__a21o_1 _3887_ (.A1(_0895_),
    .A2(_0887_),
    .B1(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__nand3_1 _3888_ (.A(_0895_),
    .B(_0887_),
    .C(_0963_),
    .Y(_0965_));
 sky130_fd_sc_hd__nand2_1 _3889_ (.A(_0964_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__or3_1 _3890_ (.A(_1354_),
    .B(_0187_),
    .C(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__o21ai_1 _3891_ (.A1(_1354_),
    .A2(_0187_),
    .B1(_0966_),
    .Y(_0968_));
 sky130_fd_sc_hd__nand2_1 _3892_ (.A(_0967_),
    .B(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__nand2b_1 _3893_ (.A_N(_0958_),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__inv_2 _3894_ (.A(_0969_),
    .Y(_0971_));
 sky130_fd_sc_hd__nand2_1 _3895_ (.A(_0958_),
    .B(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__nand2_1 _3896_ (.A(_0970_),
    .B(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__nand2_1 _3897_ (.A(_1311_),
    .B(_1496_),
    .Y(_0974_));
 sky130_fd_sc_hd__nand2_1 _3898_ (.A(_0973_),
    .B(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__nand3b_1 _3899_ (.A_N(_0974_),
    .B(_0970_),
    .C(_0972_),
    .Y(_0976_));
 sky130_fd_sc_hd__nand2_1 _3900_ (.A(_0975_),
    .B(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__nand3_1 _3901_ (.A(_0977_),
    .B(_0906_),
    .C(_0912_),
    .Y(_0978_));
 sky130_fd_sc_hd__nand2_1 _3902_ (.A(_0912_),
    .B(_0906_),
    .Y(_0979_));
 sky130_fd_sc_hd__nand3_1 _3903_ (.A(_0979_),
    .B(_0976_),
    .C(_0975_),
    .Y(_0980_));
 sky130_fd_sc_hd__nand2_1 _3904_ (.A(_0978_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__inv_2 _3905_ (.A(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__nand2_1 _3906_ (.A(_0956_),
    .B(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__nand3_1 _3907_ (.A(_0954_),
    .B(_0981_),
    .C(_0955_),
    .Y(_0984_));
 sky130_fd_sc_hd__nand2_1 _3908_ (.A(_0983_),
    .B(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__nand2_1 _3909_ (.A(_0916_),
    .B(_0567_),
    .Y(_0986_));
 sky130_fd_sc_hd__nand2_1 _3910_ (.A(_0986_),
    .B(_0915_),
    .Y(_0987_));
 sky130_fd_sc_hd__nand3_1 _3911_ (.A(_0933_),
    .B(_0985_),
    .C(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__o21ai_1 _3912_ (.A1(_0917_),
    .A2(_0571_),
    .B1(_0987_),
    .Y(_0989_));
 sky130_fd_sc_hd__inv_2 _3913_ (.A(_0985_),
    .Y(_0990_));
 sky130_fd_sc_hd__nand2_1 _3914_ (.A(_0989_),
    .B(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__nand2_1 _3915_ (.A(_0988_),
    .B(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__inv_2 _3916_ (.A(_0845_),
    .Y(_0993_));
 sky130_fd_sc_hd__nand2_1 _3917_ (.A(_0836_),
    .B(_0832_),
    .Y(_0994_));
 sky130_fd_sc_hd__nand2_1 _3918_ (.A(\datapath.MultiplierAC.PPG0.Y[11] ),
    .B(_1488_),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2_1 _3919_ (.A(\datapath.MultiplierAC.PPG0.Y[8] ),
    .B(_1494_),
    .Y(_0996_));
 sky130_fd_sc_hd__nor2_1 _3920_ (.A(_0814_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__nand2_1 _3921_ (.A(_0814_),
    .B(_0996_),
    .Y(_0998_));
 sky130_fd_sc_hd__or2b_1 _3922_ (.A(_0997_),
    .B_N(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__nand2_1 _3923_ (.A(_0822_),
    .B(_0816_),
    .Y(_1000_));
 sky130_fd_sc_hd__xor2_1 _3924_ (.A(_0999_),
    .B(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__or3_1 _3925_ (.A(_1237_),
    .B(_1657_),
    .C(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__o21ai_1 _3926_ (.A1(_1237_),
    .A2(_1657_),
    .B1(_1001_),
    .Y(_1003_));
 sky130_fd_sc_hd__nand2_1 _3927_ (.A(_1002_),
    .B(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__nand2_1 _3928_ (.A(_0830_),
    .B(_0825_),
    .Y(_1005_));
 sky130_fd_sc_hd__nand2b_1 _3929_ (.A_N(_1004_),
    .B(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__nand2b_1 _3930_ (.A_N(_1005_),
    .B(_1004_),
    .Y(_1007_));
 sky130_fd_sc_hd__nand2_1 _3931_ (.A(_1006_),
    .B(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__or2_1 _3932_ (.A(_0995_),
    .B(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__nand2_1 _3933_ (.A(_1008_),
    .B(_0995_),
    .Y(_1010_));
 sky130_fd_sc_hd__nand2_1 _3934_ (.A(_1009_),
    .B(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__inv_2 _3935_ (.A(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__nand2_1 _3936_ (.A(_0994_),
    .B(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__nand3_1 _3937_ (.A(_0836_),
    .B(_0832_),
    .C(_1011_),
    .Y(_1014_));
 sky130_fd_sc_hd__nand2_1 _3938_ (.A(_1013_),
    .B(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__nand2_1 _3939_ (.A(\datapath.MultiplierAC.PPG0.Y[12] ),
    .B(_1485_),
    .Y(_1016_));
 sky130_fd_sc_hd__xnor2_1 _3940_ (.A(_0840_),
    .B(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__xor2_1 _3941_ (.A(_0841_),
    .B(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__or3_1 _3942_ (.A(_1121_),
    .B(_1510_),
    .C(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__o21ai_1 _3943_ (.A1(_1121_),
    .A2(_1510_),
    .B1(_1018_),
    .Y(_1020_));
 sky130_fd_sc_hd__nand2_1 _3944_ (.A(_1019_),
    .B(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__nand2_1 _3945_ (.A(_1015_),
    .B(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__nand3b_1 _3946_ (.A_N(_1021_),
    .B(_1013_),
    .C(_1014_),
    .Y(_1023_));
 sky130_fd_sc_hd__nand3_1 _3947_ (.A(_0993_),
    .B(_1022_),
    .C(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__nand2_1 _3948_ (.A(_1022_),
    .B(_1023_),
    .Y(_1025_));
 sky130_fd_sc_hd__nand2_1 _3949_ (.A(_1025_),
    .B(_0845_),
    .Y(_1026_));
 sky130_fd_sc_hd__nand2_1 _3950_ (.A(_1024_),
    .B(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__nand2_1 _3951_ (.A(_1027_),
    .B(_0850_),
    .Y(_1028_));
 sky130_fd_sc_hd__inv_2 _3952_ (.A(_0850_),
    .Y(_1029_));
 sky130_fd_sc_hd__nand3_1 _3953_ (.A(_1029_),
    .B(_1024_),
    .C(_1026_),
    .Y(_1030_));
 sky130_fd_sc_hd__nand2_1 _3954_ (.A(_1028_),
    .B(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__nand2_1 _3955_ (.A(_0992_),
    .B(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__nand3b_1 _3956_ (.A_N(_1031_),
    .B(_0988_),
    .C(_0991_),
    .Y(_1033_));
 sky130_fd_sc_hd__nand2_1 _3957_ (.A(_1032_),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__inv_2 _3958_ (.A(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__nand2_1 _3959_ (.A(_0932_),
    .B(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__nand3_1 _3960_ (.A(_1034_),
    .B(_0929_),
    .C(_0921_),
    .Y(_1037_));
 sky130_fd_sc_hd__nand3_1 _3961_ (.A(_1036_),
    .B(_1037_),
    .C(_1513_),
    .Y(_1038_));
 sky130_fd_sc_hd__nand2_1 _3962_ (.A(_1504_),
    .B(_1488_),
    .Y(_1039_));
 sky130_fd_sc_hd__nand2_1 _3963_ (.A(_1502_),
    .B(_1490_),
    .Y(_1040_));
 sky130_fd_sc_hd__nand2_1 _3964_ (.A(_1498_),
    .B(_1494_),
    .Y(_1041_));
 sky130_fd_sc_hd__nand2_1 _3965_ (.A(_0746_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__o21ai_1 _3966_ (.A1(_1764_),
    .A2(_2126_),
    .B1(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__nand2_1 _3967_ (.A(_0778_),
    .B(_0747_),
    .Y(_1044_));
 sky130_fd_sc_hd__xor2_1 _3968_ (.A(_1043_),
    .B(_1044_),
    .X(_1046_));
 sky130_fd_sc_hd__or2_1 _3969_ (.A(_1040_),
    .B(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__nand2_1 _3970_ (.A(_1046_),
    .B(_1040_),
    .Y(_1048_));
 sky130_fd_sc_hd__nand2_1 _3971_ (.A(_1047_),
    .B(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__nand2_1 _3972_ (.A(_0786_),
    .B(_0781_),
    .Y(_1050_));
 sky130_fd_sc_hd__or2b_1 _3973_ (.A(_1049_),
    .B_N(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__nand2b_1 _3974_ (.A_N(_1050_),
    .B(_1049_),
    .Y(_1052_));
 sky130_fd_sc_hd__nand2_1 _3975_ (.A(_1051_),
    .B(_1052_),
    .Y(_1053_));
 sky130_fd_sc_hd__or2_1 _3976_ (.A(_1039_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__nand2_1 _3977_ (.A(_1053_),
    .B(_1039_),
    .Y(_1055_));
 sky130_fd_sc_hd__nand2_1 _3978_ (.A(_1054_),
    .B(_1055_),
    .Y(_1057_));
 sky130_fd_sc_hd__a21o_1 _3979_ (.A1(_0794_),
    .A2(_0788_),
    .B1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__nand3_1 _3980_ (.A(_1057_),
    .B(_0794_),
    .C(_0788_),
    .Y(_1059_));
 sky130_fd_sc_hd__nand2_1 _3981_ (.A(_1058_),
    .B(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__nand2_1 _3982_ (.A(\datapath.MultiplierAC.PPG0.X[14] ),
    .B(_1475_),
    .Y(_1061_));
 sky130_fd_sc_hd__nand2_1 _3983_ (.A(\datapath.MultiplierAC.PPG0.X[12] ),
    .B(_1485_),
    .Y(_1062_));
 sky130_fd_sc_hd__xnor2_1 _3984_ (.A(_0711_),
    .B(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__xor2_1 _3985_ (.A(_0712_),
    .B(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__or2_1 _3986_ (.A(_1061_),
    .B(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__nand2_1 _3987_ (.A(_1064_),
    .B(_1061_),
    .Y(_1066_));
 sky130_fd_sc_hd__nand2_1 _3988_ (.A(_1065_),
    .B(_1066_),
    .Y(_1068_));
 sky130_fd_sc_hd__nand2_1 _3989_ (.A(_1060_),
    .B(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__nand3b_1 _3990_ (.A_N(_1068_),
    .B(_1058_),
    .C(_1059_),
    .Y(_1070_));
 sky130_fd_sc_hd__nand2_1 _3991_ (.A(_1069_),
    .B(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__nand2_1 _3992_ (.A(_1071_),
    .B(_0796_),
    .Y(_1072_));
 sky130_fd_sc_hd__nand3b_1 _3993_ (.A_N(_0796_),
    .B(_1069_),
    .C(_1070_),
    .Y(_1073_));
 sky130_fd_sc_hd__inv_2 _3994_ (.A(_0800_),
    .Y(_1074_));
 sky130_fd_sc_hd__a21o_1 _3995_ (.A1(_1072_),
    .A2(_1073_),
    .B1(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__nand3_1 _3996_ (.A(_1074_),
    .B(_1073_),
    .C(_1072_),
    .Y(_1076_));
 sky130_fd_sc_hd__nand2_1 _3997_ (.A(_1075_),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__inv_2 _3998_ (.A(_0767_),
    .Y(_1079_));
 sky130_fd_sc_hd__o21a_1 _3999_ (.A1(_0660_),
    .A2(_1079_),
    .B1(_0769_),
    .X(_1080_));
 sky130_fd_sc_hd__nand3_1 _4000_ (.A(_0771_),
    .B(_0662_),
    .C(_0607_),
    .Y(_1081_));
 sky130_fd_sc_hd__nand2_1 _4001_ (.A(_1080_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__o21ai_1 _4002_ (.A1(_0651_),
    .A2(_0762_),
    .B1(_0760_),
    .Y(_1083_));
 sky130_fd_sc_hd__and3_1 _4003_ (.A(_0656_),
    .B(_0763_),
    .C(_0741_),
    .X(_1084_));
 sky130_fd_sc_hd__nor2_1 _4004_ (.A(_0746_),
    .B(_1040_),
    .Y(_1085_));
 sky130_fd_sc_hd__inv_2 _4005_ (.A(_1085_),
    .Y(_1086_));
 sky130_fd_sc_hd__nand2_1 _4006_ (.A(_0746_),
    .B(_1040_),
    .Y(_1087_));
 sky130_fd_sc_hd__and2_1 _4007_ (.A(_1086_),
    .B(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__nand2_1 _4008_ (.A(_0750_),
    .B(_0747_),
    .Y(_1090_));
 sky130_fd_sc_hd__or2_1 _4009_ (.A(_1088_),
    .B(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__nand2_1 _4010_ (.A(_1090_),
    .B(_1088_),
    .Y(_1092_));
 sky130_fd_sc_hd__nand2_1 _4011_ (.A(_1091_),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__or2_1 _4012_ (.A(_1041_),
    .B(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__nand2_1 _4013_ (.A(_1093_),
    .B(_1041_),
    .Y(_1095_));
 sky130_fd_sc_hd__nand2_1 _4014_ (.A(_1094_),
    .B(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__and2_1 _4015_ (.A(_0756_),
    .B(_0753_),
    .X(_1097_));
 sky130_fd_sc_hd__or2_1 _4016_ (.A(_1096_),
    .B(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__nand2_1 _4017_ (.A(_1097_),
    .B(_1096_),
    .Y(_1099_));
 sky130_fd_sc_hd__nand2_1 _4018_ (.A(_1098_),
    .B(_1099_),
    .Y(_1101_));
 sky130_fd_sc_hd__or2_1 _4019_ (.A(_0460_),
    .B(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__nand2_1 _4020_ (.A(_1101_),
    .B(_0460_),
    .Y(_1103_));
 sky130_fd_sc_hd__nand2_1 _4021_ (.A(_1102_),
    .B(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__o21bai_1 _4022_ (.A1(_1083_),
    .A2(_1084_),
    .B1_N(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__nor2_1 _4023_ (.A(_1083_),
    .B(_1084_),
    .Y(_1106_));
 sky130_fd_sc_hd__nand2_1 _4024_ (.A(_1106_),
    .B(_1104_),
    .Y(_1107_));
 sky130_fd_sc_hd__nand2_1 _4025_ (.A(_1105_),
    .B(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__nand2_1 _4026_ (.A(_0738_),
    .B(_0735_),
    .Y(_1109_));
 sky130_fd_sc_hd__or2_1 _4027_ (.A(_0711_),
    .B(_1061_),
    .X(_1110_));
 sky130_fd_sc_hd__nand2_1 _4028_ (.A(_0711_),
    .B(_1061_),
    .Y(_1111_));
 sky130_fd_sc_hd__nand2_1 _4029_ (.A(_1110_),
    .B(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__nand2_1 _4030_ (.A(_0723_),
    .B(_0713_),
    .Y(_1113_));
 sky130_fd_sc_hd__xor2_1 _4031_ (.A(_1112_),
    .B(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__or2_1 _4032_ (.A(_1062_),
    .B(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__nand2_1 _4033_ (.A(_1114_),
    .B(_1062_),
    .Y(_1116_));
 sky130_fd_sc_hd__nand2_1 _4034_ (.A(_1115_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__inv_2 _4035_ (.A(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__o21ai_1 _4036_ (.A1(_0728_),
    .A2(_0627_),
    .B1(_0727_),
    .Y(_1119_));
 sky130_fd_sc_hd__nand3_1 _4037_ (.A(_0626_),
    .B(_0627_),
    .C(_0729_),
    .Y(_1120_));
 sky130_fd_sc_hd__nor2_1 _4038_ (.A(_0612_),
    .B(_1120_),
    .Y(_1122_));
 sky130_fd_sc_hd__nor2_1 _4039_ (.A(_1119_),
    .B(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__inv_2 _4040_ (.A(_1120_),
    .Y(_1124_));
 sky130_fd_sc_hd__nand3_1 _4041_ (.A(_1124_),
    .B(_0268_),
    .C(_0609_),
    .Y(_1125_));
 sky130_fd_sc_hd__nand2_1 _4042_ (.A(_1123_),
    .B(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__or2_1 _4043_ (.A(_1118_),
    .B(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__nand2_1 _4044_ (.A(_1126_),
    .B(_1118_),
    .Y(_1128_));
 sky130_fd_sc_hd__nand2_1 _4045_ (.A(_1127_),
    .B(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__nand2_1 _4046_ (.A(_1129_),
    .B(_1039_),
    .Y(_1130_));
 sky130_fd_sc_hd__nand3b_1 _4047_ (.A_N(_1039_),
    .B(_1127_),
    .C(_1128_),
    .Y(_1131_));
 sky130_fd_sc_hd__nand2_1 _4048_ (.A(_1130_),
    .B(_1131_),
    .Y(_1133_));
 sky130_fd_sc_hd__inv_2 _4049_ (.A(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__nand2_1 _4050_ (.A(_1109_),
    .B(_1134_),
    .Y(_1135_));
 sky130_fd_sc_hd__nand3_1 _4051_ (.A(_1133_),
    .B(_0738_),
    .C(_0735_),
    .Y(_1136_));
 sky130_fd_sc_hd__nand3b_1 _4052_ (.A_N(_1108_),
    .B(_1135_),
    .C(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__nand2_1 _4053_ (.A(_1135_),
    .B(_1136_),
    .Y(_1138_));
 sky130_fd_sc_hd__nand2_1 _4054_ (.A(_1138_),
    .B(_1108_),
    .Y(_1139_));
 sky130_fd_sc_hd__nand2_1 _4055_ (.A(_1137_),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__inv_2 _4056_ (.A(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__nand2_1 _4057_ (.A(_1082_),
    .B(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__nand3_1 _4058_ (.A(_1140_),
    .B(_1080_),
    .C(_1081_),
    .Y(_1143_));
 sky130_fd_sc_hd__nand3b_1 _4059_ (.A_N(_1077_),
    .B(_1142_),
    .C(_1143_),
    .Y(_1144_));
 sky130_fd_sc_hd__nand2_1 _4060_ (.A(_1142_),
    .B(_1143_),
    .Y(_1145_));
 sky130_fd_sc_hd__nand2_1 _4061_ (.A(_1145_),
    .B(_1077_),
    .Y(_1146_));
 sky130_fd_sc_hd__nand2_1 _4062_ (.A(_1144_),
    .B(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__inv_2 _4063_ (.A(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__nand2_1 _4064_ (.A(_0809_),
    .B(_0805_),
    .Y(_1149_));
 sky130_fd_sc_hd__or2_1 _4065_ (.A(_1148_),
    .B(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__nand2_1 _4066_ (.A(_1149_),
    .B(_1148_),
    .Y(_1151_));
 sky130_fd_sc_hd__nand3_1 _4067_ (.A(_1150_),
    .B(_1538_),
    .C(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__nand2_1 _4068_ (.A(_1038_),
    .B(_1152_),
    .Y(_1154_));
 sky130_fd_sc_hd__nand2_1 _4069_ (.A(_1154_),
    .B(_1517_),
    .Y(_1155_));
 sky130_fd_sc_hd__nand2_1 _4070_ (.A(_1518_),
    .B(\datapath.MultiplierAC.PPG0.X[13] ),
    .Y(_1156_));
 sky130_fd_sc_hd__a21oi_1 _4071_ (.A1(_1155_),
    .A2(_1156_),
    .B1(_1545_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand2_1 _4072_ (.A(_1151_),
    .B(_1144_),
    .Y(_1157_));
 sky130_fd_sc_hd__nand2_1 _4073_ (.A(_1076_),
    .B(_1073_),
    .Y(_1158_));
 sky130_fd_sc_hd__nand2_1 _4074_ (.A(_1504_),
    .B(_1490_),
    .Y(_1159_));
 sky130_fd_sc_hd__nand2_1 _4075_ (.A(_1502_),
    .B(_1492_),
    .Y(_1160_));
 sky130_fd_sc_hd__nand2_1 _4076_ (.A(_1500_),
    .B(_1494_),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _4077_ (.A(_2059_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__o21a_1 _4078_ (.A1(_1929_),
    .A2(_2126_),
    .B1(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__nor2_1 _4079_ (.A(_1764_),
    .B(_2126_),
    .Y(_1164_));
 sky130_fd_sc_hd__o21ai_1 _4080_ (.A1(_1164_),
    .A2(_1044_),
    .B1(_1042_),
    .Y(_1165_));
 sky130_fd_sc_hd__xor2_1 _4081_ (.A(_1163_),
    .B(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__xnor2_1 _4082_ (.A(_1160_),
    .B(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__nand2_1 _4083_ (.A(_1051_),
    .B(_1047_),
    .Y(_1168_));
 sky130_fd_sc_hd__xor2_1 _4084_ (.A(_1167_),
    .B(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__xor2_1 _4085_ (.A(_1159_),
    .B(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__nand3b_1 _4086_ (.A_N(_1170_),
    .B(_1054_),
    .C(_1058_),
    .Y(_1171_));
 sky130_fd_sc_hd__nand2_1 _4087_ (.A(_1058_),
    .B(_1054_),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_1 _4088_ (.A(_1172_),
    .B(_1170_),
    .Y(_1174_));
 sky130_fd_sc_hd__nand2_1 _4089_ (.A(_1171_),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__nand2_1 _4090_ (.A(\datapath.MultiplierAC.PPG0.X[15] ),
    .B(_1475_),
    .Y(_1176_));
 sky130_fd_sc_hd__nand2_1 _4091_ (.A(\datapath.MultiplierAC.PPG0.X[14] ),
    .B(_1482_),
    .Y(_1177_));
 sky130_fd_sc_hd__a21oi_1 _4092_ (.A1(_0615_),
    .A2(_1062_),
    .B1(_0711_),
    .Y(_1178_));
 sky130_fd_sc_hd__nand2_1 _4093_ (.A(\datapath.MultiplierAC.PPG0.X[13] ),
    .B(_1485_),
    .Y(_1179_));
 sky130_fd_sc_hd__nand2_1 _4094_ (.A(\datapath.MultiplierAC.PPG0.X[12] ),
    .B(_1488_),
    .Y(_1180_));
 sky130_fd_sc_hd__xnor2_1 _4095_ (.A(_1179_),
    .B(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__xor2_1 _4096_ (.A(_1178_),
    .B(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__xnor2_1 _4097_ (.A(_1177_),
    .B(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__xnor2_1 _4098_ (.A(_1065_),
    .B(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__xnor2_1 _4099_ (.A(_1176_),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__nand2_1 _4100_ (.A(_1175_),
    .B(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__nand3b_1 _4101_ (.A_N(_1185_),
    .B(_1171_),
    .C(_1174_),
    .Y(_1187_));
 sky130_fd_sc_hd__nand3b_1 _4102_ (.A_N(_1070_),
    .B(_1186_),
    .C(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__nand2_1 _4103_ (.A(_1186_),
    .B(_1187_),
    .Y(_1189_));
 sky130_fd_sc_hd__nand2_1 _4104_ (.A(_1189_),
    .B(_1070_),
    .Y(_1190_));
 sky130_fd_sc_hd__nand3_1 _4105_ (.A(_1158_),
    .B(_1188_),
    .C(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__inv_2 _4106_ (.A(_1158_),
    .Y(_1192_));
 sky130_fd_sc_hd__nand2_1 _4107_ (.A(_1190_),
    .B(_1188_),
    .Y(_1193_));
 sky130_fd_sc_hd__nand2_1 _4108_ (.A(_1192_),
    .B(_1193_),
    .Y(_1195_));
 sky130_fd_sc_hd__nand2_1 _4109_ (.A(_1191_),
    .B(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__nand2_1 _4110_ (.A(_1142_),
    .B(_1137_),
    .Y(_1197_));
 sky130_fd_sc_hd__nand2_1 _4111_ (.A(_1135_),
    .B(_1131_),
    .Y(_1198_));
 sky130_fd_sc_hd__xor2_1 _4112_ (.A(_1177_),
    .B(_1176_),
    .X(_1199_));
 sky130_fd_sc_hd__o211a_1 _4113_ (.A1(_1112_),
    .A2(_0723_),
    .B1(_0713_),
    .C1(_1110_),
    .X(_1200_));
 sky130_fd_sc_hd__xor2_1 _4114_ (.A(_1199_),
    .B(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__xnor2_1 _4115_ (.A(_1179_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__nand2_1 _4116_ (.A(_1128_),
    .B(_1115_),
    .Y(_1203_));
 sky130_fd_sc_hd__xor2_1 _4117_ (.A(_1202_),
    .B(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__or2_1 _4118_ (.A(_1180_),
    .B(_1204_),
    .X(_1206_));
 sky130_fd_sc_hd__nand2_1 _4119_ (.A(_1204_),
    .B(_1180_),
    .Y(_1207_));
 sky130_fd_sc_hd__nand3_1 _4120_ (.A(_1198_),
    .B(_1206_),
    .C(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__inv_2 _4121_ (.A(_1180_),
    .Y(_1209_));
 sky130_fd_sc_hd__xor2_1 _4122_ (.A(_1209_),
    .B(_1204_),
    .X(_1210_));
 sky130_fd_sc_hd__nand3_1 _4123_ (.A(_1210_),
    .B(_1131_),
    .C(_1135_),
    .Y(_1211_));
 sky130_fd_sc_hd__nand2_1 _4124_ (.A(_1208_),
    .B(_1211_),
    .Y(_1212_));
 sky130_fd_sc_hd__nand2_1 _4125_ (.A(_1105_),
    .B(_1102_),
    .Y(_1213_));
 sky130_fd_sc_hd__xnor2_1 _4126_ (.A(_1160_),
    .B(_1159_),
    .Y(_1214_));
 sky130_fd_sc_hd__nand2_1 _4127_ (.A(_1092_),
    .B(_1086_),
    .Y(_1215_));
 sky130_fd_sc_hd__xor2_1 _4128_ (.A(_1214_),
    .B(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__xnor2_1 _4129_ (.A(_1161_),
    .B(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__nand2_1 _4130_ (.A(_1098_),
    .B(_1094_),
    .Y(_1218_));
 sky130_fd_sc_hd__xor2_1 _4131_ (.A(_1217_),
    .B(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__xor2_1 _4132_ (.A(_2060_),
    .B(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__inv_2 _4133_ (.A(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__nand2_1 _4134_ (.A(_1213_),
    .B(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__nand3_1 _4135_ (.A(_1105_),
    .B(_1102_),
    .C(_1220_),
    .Y(_1223_));
 sky130_fd_sc_hd__nand2_1 _4136_ (.A(_1222_),
    .B(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__nand2_1 _4137_ (.A(_1212_),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__inv_2 _4138_ (.A(_1224_),
    .Y(_1227_));
 sky130_fd_sc_hd__nand3_1 _4139_ (.A(_1227_),
    .B(_1208_),
    .C(_1211_),
    .Y(_1228_));
 sky130_fd_sc_hd__nand2_1 _4140_ (.A(_1225_),
    .B(_1228_),
    .Y(_1229_));
 sky130_fd_sc_hd__inv_2 _4141_ (.A(_1229_),
    .Y(_1230_));
 sky130_fd_sc_hd__nand2_1 _4142_ (.A(_1197_),
    .B(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__nand3_1 _4143_ (.A(_1229_),
    .B(_1142_),
    .C(_1137_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand3b_1 _4144_ (.A_N(_1196_),
    .B(_1231_),
    .C(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__nand2_1 _4145_ (.A(_1231_),
    .B(_1232_),
    .Y(_1234_));
 sky130_fd_sc_hd__nand2_1 _4146_ (.A(_1234_),
    .B(_1196_),
    .Y(_1235_));
 sky130_fd_sc_hd__nand2_1 _4147_ (.A(_1233_),
    .B(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__inv_2 _4148_ (.A(_1236_),
    .Y(_1238_));
 sky130_fd_sc_hd__nand2_1 _4149_ (.A(_1157_),
    .B(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__nand3_1 _4150_ (.A(_1151_),
    .B(_1236_),
    .C(_1144_),
    .Y(_1240_));
 sky130_fd_sc_hd__nand3_1 _4151_ (.A(_1239_),
    .B(_1538_),
    .C(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__nand2_1 _4152_ (.A(_1241_),
    .B(_1517_),
    .Y(_1242_));
 sky130_fd_sc_hd__inv_2 _4153_ (.A(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__nand2_1 _4154_ (.A(_1036_),
    .B(_1033_),
    .Y(_1244_));
 sky130_fd_sc_hd__nand2_1 _4155_ (.A(_0991_),
    .B(_0983_),
    .Y(_1245_));
 sky130_fd_sc_hd__nor2_1 _4156_ (.A(_0879_),
    .B(_0952_),
    .Y(_1246_));
 sky130_fd_sc_hd__nand2_1 _4157_ (.A(_1246_),
    .B(_0855_),
    .Y(_1247_));
 sky130_fd_sc_hd__inv_2 _4158_ (.A(_0875_),
    .Y(_1249_));
 sky130_fd_sc_hd__a21boi_1 _4159_ (.A1(_0950_),
    .A2(_1249_),
    .B1_N(_0951_),
    .Y(_1250_));
 sky130_fd_sc_hd__nand2_1 _4160_ (.A(_1247_),
    .B(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__nand2_1 _4161_ (.A(_1435_),
    .B(\datapath.MultiplierAC.PPG0.X[12] ),
    .Y(_1252_));
 sky130_fd_sc_hd__nand2_1 _4162_ (.A(_0947_),
    .B(_0941_),
    .Y(_1253_));
 sky130_fd_sc_hd__nand2_1 _4163_ (.A(_1448_),
    .B(\datapath.MultiplierAC.PPG0.X[13] ),
    .Y(_1254_));
 sky130_fd_sc_hd__nand2_1 _4164_ (.A(_1463_),
    .B(\datapath.MultiplierAC.PPG0.X[15] ),
    .Y(_1255_));
 sky130_fd_sc_hd__a22o_1 _4165_ (.A1(_1463_),
    .A2(\datapath.MultiplierAC.PPG0.X[14] ),
    .B1(_1466_),
    .B2(\datapath.MultiplierAC.PPG0.X[15] ),
    .X(_1256_));
 sky130_fd_sc_hd__o21ai_1 _4166_ (.A1(_0937_),
    .A2(_1255_),
    .B1(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__a21o_1 _4167_ (.A1(_0516_),
    .A2(_0937_),
    .B1(_0857_),
    .X(_1258_));
 sky130_fd_sc_hd__o21ai_1 _4168_ (.A1(_0938_),
    .A2(_0865_),
    .B1(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__xor2_1 _4169_ (.A(_1257_),
    .B(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__xnor2_1 _4170_ (.A(_1254_),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__or2b_1 _4171_ (.A(_1253_),
    .B_N(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__a21o_1 _4172_ (.A1(_0947_),
    .A2(_0941_),
    .B1(_1261_),
    .X(_1263_));
 sky130_fd_sc_hd__nand3b_1 _4173_ (.A_N(_1252_),
    .B(_1262_),
    .C(_1263_),
    .Y(_1264_));
 sky130_fd_sc_hd__or2_1 _4174_ (.A(_1261_),
    .B(_1253_),
    .X(_1265_));
 sky130_fd_sc_hd__nand2_1 _4175_ (.A(_1253_),
    .B(_1261_),
    .Y(_1266_));
 sky130_fd_sc_hd__nand3_1 _4176_ (.A(_1265_),
    .B(_1252_),
    .C(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__nand2_1 _4177_ (.A(_1264_),
    .B(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__inv_2 _4178_ (.A(_1268_),
    .Y(_1270_));
 sky130_fd_sc_hd__nand2_1 _4179_ (.A(_1251_),
    .B(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__nand3_1 _4180_ (.A(_1247_),
    .B(_1268_),
    .C(_1250_),
    .Y(_1272_));
 sky130_fd_sc_hd__nand2_1 _4181_ (.A(_1271_),
    .B(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__nand2_1 _4182_ (.A(_0980_),
    .B(_0976_),
    .Y(_1274_));
 sky130_fd_sc_hd__nand2_1 _4183_ (.A(_0972_),
    .B(_0967_),
    .Y(_1275_));
 sky130_fd_sc_hd__nand2_1 _4184_ (.A(_1343_),
    .B(_1500_),
    .Y(_1276_));
 sky130_fd_sc_hd__inv_2 _4185_ (.A(_1276_),
    .Y(_1277_));
 sky130_fd_sc_hd__nand2_1 _4186_ (.A(_1379_),
    .B(_1504_),
    .Y(_1278_));
 sky130_fd_sc_hd__a22o_1 _4187_ (.A1(_1379_),
    .A2(_1502_),
    .B1(_1411_),
    .B2(_1504_),
    .X(_1279_));
 sky130_fd_sc_hd__o21a_1 _4188_ (.A1(_0959_),
    .A2(_1278_),
    .B1(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__nand2_1 _4189_ (.A(_0964_),
    .B(_0961_),
    .Y(_1281_));
 sky130_fd_sc_hd__xnor2_1 _4190_ (.A(_1280_),
    .B(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__xor2_1 _4191_ (.A(_1277_),
    .B(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__inv_2 _4192_ (.A(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__nand2_1 _4193_ (.A(_1275_),
    .B(_1284_),
    .Y(_1285_));
 sky130_fd_sc_hd__nand3_1 _4194_ (.A(_0972_),
    .B(_0967_),
    .C(_1283_),
    .Y(_1286_));
 sky130_fd_sc_hd__nand2_1 _4195_ (.A(_1285_),
    .B(_1286_),
    .Y(_1287_));
 sky130_fd_sc_hd__nand2_1 _4196_ (.A(_1311_),
    .B(_1498_),
    .Y(_1288_));
 sky130_fd_sc_hd__nand2_1 _4197_ (.A(_1287_),
    .B(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__inv_2 _4198_ (.A(_1288_),
    .Y(_1291_));
 sky130_fd_sc_hd__nand3_1 _4199_ (.A(_1285_),
    .B(_1291_),
    .C(_1286_),
    .Y(_1292_));
 sky130_fd_sc_hd__nand2_1 _4200_ (.A(_1289_),
    .B(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__inv_2 _4201_ (.A(_1293_),
    .Y(_1294_));
 sky130_fd_sc_hd__nand2_1 _4202_ (.A(_1274_),
    .B(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__nand3_1 _4203_ (.A(_0980_),
    .B(_1293_),
    .C(_0976_),
    .Y(_1296_));
 sky130_fd_sc_hd__nand2_1 _4204_ (.A(_1295_),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__nand2_1 _4205_ (.A(_1273_),
    .B(_1297_),
    .Y(_1298_));
 sky130_fd_sc_hd__inv_2 _4206_ (.A(_1297_),
    .Y(_1299_));
 sky130_fd_sc_hd__nand3_1 _4207_ (.A(_1299_),
    .B(_1271_),
    .C(_1272_),
    .Y(_1300_));
 sky130_fd_sc_hd__nand2_1 _4208_ (.A(_1298_),
    .B(_1300_),
    .Y(_1301_));
 sky130_fd_sc_hd__nand2_1 _4209_ (.A(_1245_),
    .B(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__nand2_1 _4210_ (.A(_1273_),
    .B(_1299_),
    .Y(_1303_));
 sky130_fd_sc_hd__nand3_1 _4211_ (.A(_1271_),
    .B(_1272_),
    .C(_1297_),
    .Y(_1304_));
 sky130_fd_sc_hd__nand2_1 _4212_ (.A(_1303_),
    .B(_1304_),
    .Y(_1305_));
 sky130_fd_sc_hd__nand3_1 _4213_ (.A(_0991_),
    .B(_1305_),
    .C(_0983_),
    .Y(_1306_));
 sky130_fd_sc_hd__nand2_1 _4214_ (.A(_1302_),
    .B(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__nand2_1 _4215_ (.A(\datapath.MultiplierAC.PPG0.Y[11] ),
    .B(_1490_),
    .Y(_1308_));
 sky130_fd_sc_hd__nand2_1 _4216_ (.A(\datapath.MultiplierAC.PPG0.Y[10] ),
    .B(_1492_),
    .Y(_1309_));
 sky130_fd_sc_hd__nand2_1 _4217_ (.A(\datapath.MultiplierAC.PPG0.Y[9] ),
    .B(_1496_),
    .Y(_1310_));
 sky130_fd_sc_hd__a22o_1 _4218_ (.A1(\datapath.MultiplierAC.PPG0.Y[9] ),
    .A2(_1494_),
    .B1(\datapath.MultiplierAC.PPG0.Y[8] ),
    .B2(_1496_),
    .X(_1312_));
 sky130_fd_sc_hd__o21ai_1 _4219_ (.A1(_0996_),
    .A2(_1310_),
    .B1(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__nor2_1 _4220_ (.A(_0999_),
    .B(_0817_),
    .Y(_1314_));
 sky130_fd_sc_hd__a211o_1 _4221_ (.A1(_0820_),
    .A2(_1314_),
    .B1(_0815_),
    .C1(_0997_),
    .X(_1315_));
 sky130_fd_sc_hd__xor2_1 _4222_ (.A(_1313_),
    .B(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__xor2_1 _4223_ (.A(_1309_),
    .B(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__nand2_1 _4224_ (.A(_1006_),
    .B(_1002_),
    .Y(_1318_));
 sky130_fd_sc_hd__xor2_1 _4225_ (.A(_1317_),
    .B(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__xnor2_1 _4226_ (.A(_1308_),
    .B(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__nand3b_1 _4227_ (.A_N(_1320_),
    .B(_1009_),
    .C(_1013_),
    .Y(_1321_));
 sky130_fd_sc_hd__nand2_1 _4228_ (.A(_1013_),
    .B(_1009_),
    .Y(_1323_));
 sky130_fd_sc_hd__nand2_1 _4229_ (.A(_1323_),
    .B(_1320_),
    .Y(_1324_));
 sky130_fd_sc_hd__nand2_1 _4230_ (.A(_1321_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_1 _4231_ (.A(\datapath.MultiplierAC.PPG0.Y[15] ),
    .B(_1475_),
    .Y(_1326_));
 sky130_fd_sc_hd__nand2_1 _4232_ (.A(\datapath.MultiplierAC.PPG0.Y[14] ),
    .B(_1482_),
    .Y(_1327_));
 sky130_fd_sc_hd__a21oi_1 _4233_ (.A1(_0574_),
    .A2(_1016_),
    .B1(_0840_),
    .Y(_1328_));
 sky130_fd_sc_hd__nand2_1 _4234_ (.A(\datapath.MultiplierAC.PPG0.Y[13] ),
    .B(_1488_),
    .Y(_1329_));
 sky130_fd_sc_hd__a22o_1 _4235_ (.A1(\datapath.MultiplierAC.PPG0.Y[13] ),
    .A2(_1485_),
    .B1(\datapath.MultiplierAC.PPG0.Y[12] ),
    .B2(_1488_),
    .X(_1330_));
 sky130_fd_sc_hd__o21ai_1 _4236_ (.A1(_1016_),
    .A2(_1329_),
    .B1(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__xor2_1 _4237_ (.A(_1328_),
    .B(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__xnor2_1 _4238_ (.A(_1327_),
    .B(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__xnor2_1 _4239_ (.A(_1019_),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__xnor2_1 _4240_ (.A(_1326_),
    .B(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__nand2_1 _4241_ (.A(_1325_),
    .B(_1335_),
    .Y(_1336_));
 sky130_fd_sc_hd__nand3b_1 _4242_ (.A_N(_1335_),
    .B(_1321_),
    .C(_1324_),
    .Y(_1337_));
 sky130_fd_sc_hd__nand2_1 _4243_ (.A(_1336_),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__nand2_1 _4244_ (.A(_1338_),
    .B(_1023_),
    .Y(_1339_));
 sky130_fd_sc_hd__nand3b_1 _4245_ (.A_N(_1023_),
    .B(_1336_),
    .C(_1337_),
    .Y(_1340_));
 sky130_fd_sc_hd__nand2_1 _4246_ (.A(_1339_),
    .B(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__nand2_1 _4247_ (.A(_1030_),
    .B(_1024_),
    .Y(_1342_));
 sky130_fd_sc_hd__inv_2 _4248_ (.A(_1342_),
    .Y(_1344_));
 sky130_fd_sc_hd__nand2_1 _4249_ (.A(_1341_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__nand3_1 _4250_ (.A(_1342_),
    .B(_1339_),
    .C(_1340_),
    .Y(_1346_));
 sky130_fd_sc_hd__nand2_1 _4251_ (.A(_1345_),
    .B(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__inv_2 _4252_ (.A(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__nand2_1 _4253_ (.A(_1307_),
    .B(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__nand3_1 _4254_ (.A(_1302_),
    .B(_1306_),
    .C(_1347_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand2_1 _4255_ (.A(_1349_),
    .B(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__inv_2 _4256_ (.A(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__nand2_1 _4257_ (.A(_1244_),
    .B(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__nand3_1 _4258_ (.A(_1036_),
    .B(_1351_),
    .C(_1033_),
    .Y(_1355_));
 sky130_fd_sc_hd__nand3_1 _4259_ (.A(_1353_),
    .B(_1513_),
    .C(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__o21ai_1 _4260_ (.A1(_1517_),
    .A2(\datapath.MultiplierAC.PPG0.X[14] ),
    .B1(_1067_),
    .Y(_1357_));
 sky130_fd_sc_hd__a21oi_1 _4261_ (.A1(_1243_),
    .A2(_1356_),
    .B1(_1357_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _4262_ (.A(\control_unit.state[2] ),
    .Y(_1358_));
 sky130_fd_sc_hd__inv_2 _4263_ (.A(\control_unit.state[1] ),
    .Y(_1359_));
 sky130_fd_sc_hd__and3_1 _4264_ (.A(_1358_),
    .B(_1359_),
    .C(\control_unit.state[0] ),
    .X(_1360_));
 sky130_fd_sc_hd__nor2_1 _4265_ (.A(\control_unit.state[2] ),
    .B(_1359_),
    .Y(_1361_));
 sky130_fd_sc_hd__nor2_1 _4266_ (.A(\control_unit.state[1] ),
    .B(_1358_),
    .Y(_1362_));
 sky130_fd_sc_hd__nor2_1 _4267_ (.A(_1361_),
    .B(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__inv_2 _4268_ (.A(_1363_),
    .Y(_1365_));
 sky130_fd_sc_hd__nor2_2 _4269_ (.A(_1360_),
    .B(_1365_),
    .Y(_1366_));
 sky130_fd_sc_hd__inv_2 _4270_ (.A(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__inv_2 _4271_ (.A(_1361_),
    .Y(_1368_));
 sky130_fd_sc_hd__nor2_1 _4272_ (.A(\control_unit.state[0] ),
    .B(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__nand2_1 _4273_ (.A(_1478_),
    .B(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__o21ai_1 _4274_ (.A1(_1537_),
    .A2(_1367_),
    .B1(_1370_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _4275_ (.A(_1362_),
    .Y(_1371_));
 sky130_fd_sc_hd__nor2_1 _4276_ (.A(\control_unit.state[0] ),
    .B(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__nand2_1 _4277_ (.A(_1372_),
    .B(\control_unit.regBk ),
    .Y(_1373_));
 sky130_fd_sc_hd__inv_2 _4278_ (.A(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__a21o_1 _4279_ (.A1(_1366_),
    .A2(\control_unit.S_C[1] ),
    .B1(_1374_),
    .X(_0033_));
 sky130_fd_sc_hd__a21o_1 _4280_ (.A1(_1366_),
    .A2(\control_unit.S_Coun ),
    .B1(_1369_),
    .X(_0034_));
 sky130_fd_sc_hd__a32o_1 _4281_ (.A1(_1370_),
    .A2(_1373_),
    .A3(_1365_),
    .B1(_1518_),
    .B2(_1366_),
    .X(_1375_));
 sky130_fd_sc_hd__clkinv_2 _4282_ (.A(_1375_),
    .Y(_0035_));
 sky130_fd_sc_hd__buf_6 _4283_ (.A(\control_unit.ShiftB ),
    .X(_1376_));
 sky130_fd_sc_hd__a21o_1 _4284_ (.A1(_1366_),
    .A2(_1376_),
    .B1(_1372_),
    .X(_0036_));
 sky130_fd_sc_hd__a22o_1 _4285_ (.A1(net34),
    .A2(_1360_),
    .B1(_1366_),
    .B2(_1089_),
    .X(_0037_));
 sky130_fd_sc_hd__nand2_1 _4286_ (.A(_1363_),
    .B(net34),
    .Y(_1377_));
 sky130_fd_sc_hd__nand2_1 _4287_ (.A(_1367_),
    .B(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__o22a_1 _4288_ (.A1(\control_unit.LoadCoun ),
    .A2(_1367_),
    .B1(_1369_),
    .B2(_1378_),
    .X(_0038_));
 sky130_fd_sc_hd__inv_2 _4289_ (.A(\control_unit.state[0] ),
    .Y(_1380_));
 sky130_fd_sc_hd__nor2_1 _4290_ (.A(_1380_),
    .B(_1368_),
    .Y(_1381_));
 sky130_fd_sc_hd__a21o_1 _4291_ (.A1(\control_unit.regBk ),
    .A2(_1380_),
    .B1(_1371_),
    .X(_1382_));
 sky130_fd_sc_hd__a32o_1 _4292_ (.A1(_1367_),
    .A2(_1382_),
    .A3(_1377_),
    .B1(\control_unit.state[1] ),
    .B2(\control_unit.state[0] ),
    .X(_1383_));
 sky130_fd_sc_hd__and2b_1 _4293_ (.A_N(_1381_),
    .B(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__clkbuf_1 _4294_ (.A(_1384_),
    .X(_0039_));
 sky130_fd_sc_hd__a31o_1 _4295_ (.A1(_1382_),
    .A2(_1370_),
    .A3(_1377_),
    .B1(_1366_),
    .X(_1385_));
 sky130_fd_sc_hd__nand2_1 _4296_ (.A(\control_unit.state[2] ),
    .B(\control_unit.state[1] ),
    .Y(_1386_));
 sky130_fd_sc_hd__nand2_1 _4297_ (.A(_1385_),
    .B(_1386_),
    .Y(_0040_));
 sky130_fd_sc_hd__or3b_1 _4298_ (.A(_1381_),
    .B(_1374_),
    .C_N(_1386_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _4299_ (.A(_1388_),
    .X(_0041_));
 sky130_fd_sc_hd__and2b_1 _4300_ (.A_N(_1360_),
    .B(net51),
    .X(_1389_));
 sky130_fd_sc_hd__a21o_1 _4301_ (.A1(_1479_),
    .A2(_1369_),
    .B1(_1389_),
    .X(_0042_));
 sky130_fd_sc_hd__nor2_8 _4302_ (.A(\control_unit.LoadA ),
    .B(_1376_),
    .Y(_1390_));
 sky130_fd_sc_hd__a22o_1 _4303_ (.A1(\control_unit.LoadA ),
    .A2(net17),
    .B1(_1390_),
    .B2(\datapath.RegB[0] ),
    .X(_1391_));
 sky130_fd_sc_hd__and2_1 _4304_ (.A(_1391_),
    .B(_1067_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _4305_ (.A(_1392_),
    .X(_0043_));
 sky130_fd_sc_hd__a21o_1 _4306_ (.A1(\datapath.RegB[0] ),
    .A2(_1376_),
    .B1(_1089_),
    .X(_1393_));
 sky130_fd_sc_hd__o21ai_1 _4307_ (.A1(_1226_),
    .A2(net24),
    .B1(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__nand2_1 _4308_ (.A(_1390_),
    .B(\datapath.RegB[1] ),
    .Y(_1396_));
 sky130_fd_sc_hd__a21oi_1 _4309_ (.A1(_1394_),
    .A2(_1396_),
    .B1(_1545_),
    .Y(_0044_));
 sky130_fd_sc_hd__a21o_1 _4310_ (.A1(\datapath.RegB[1] ),
    .A2(_1376_),
    .B1(_1089_),
    .X(_1397_));
 sky130_fd_sc_hd__o21ai_1 _4311_ (.A1(_1226_),
    .A2(net25),
    .B1(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__nand2_1 _4312_ (.A(_1390_),
    .B(\datapath.RegB[2] ),
    .Y(_1399_));
 sky130_fd_sc_hd__a21oi_1 _4313_ (.A1(_1398_),
    .A2(_1399_),
    .B1(_1545_),
    .Y(_0045_));
 sky130_fd_sc_hd__a21o_1 _4314_ (.A1(\datapath.RegB[2] ),
    .A2(_1376_),
    .B1(_1089_),
    .X(_1400_));
 sky130_fd_sc_hd__o21ai_1 _4315_ (.A1(_1226_),
    .A2(net26),
    .B1(_1400_),
    .Y(_1401_));
 sky130_fd_sc_hd__nand2_1 _4316_ (.A(_1390_),
    .B(\datapath.RegB[3] ),
    .Y(_1402_));
 sky130_fd_sc_hd__a21oi_1 _4317_ (.A1(_1401_),
    .A2(_1402_),
    .B1(_1545_),
    .Y(_0046_));
 sky130_fd_sc_hd__a21o_1 _4318_ (.A1(\datapath.RegB[3] ),
    .A2(_1376_),
    .B1(_1089_),
    .X(_1403_));
 sky130_fd_sc_hd__o21ai_1 _4319_ (.A1(_1226_),
    .A2(net27),
    .B1(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__nand2_1 _4320_ (.A(_1390_),
    .B(\datapath.RegB[4] ),
    .Y(_1405_));
 sky130_fd_sc_hd__a21oi_1 _4321_ (.A1(_1404_),
    .A2(_1405_),
    .B1(_1545_),
    .Y(_0047_));
 sky130_fd_sc_hd__a21o_1 _4322_ (.A1(\datapath.RegB[4] ),
    .A2(_1376_),
    .B1(_1089_),
    .X(_1406_));
 sky130_fd_sc_hd__o21ai_1 _4323_ (.A1(_1226_),
    .A2(net28),
    .B1(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__nand2_1 _4324_ (.A(_1390_),
    .B(\datapath.RegB[5] ),
    .Y(_1408_));
 sky130_fd_sc_hd__a21oi_1 _4325_ (.A1(_1407_),
    .A2(_1408_),
    .B1(_1545_),
    .Y(_0048_));
 sky130_fd_sc_hd__a21o_1 _4326_ (.A1(\datapath.RegB[5] ),
    .A2(_1376_),
    .B1(_1089_),
    .X(_1409_));
 sky130_fd_sc_hd__o21ai_1 _4327_ (.A1(_1226_),
    .A2(net29),
    .B1(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hd__nand2_1 _4328_ (.A(_1390_),
    .B(\datapath.RegB[6] ),
    .Y(_1412_));
 sky130_fd_sc_hd__a21oi_1 _4329_ (.A1(_1410_),
    .A2(_1412_),
    .B1(_1545_),
    .Y(_0049_));
 sky130_fd_sc_hd__a21o_1 _4330_ (.A1(\datapath.RegB[6] ),
    .A2(_1376_),
    .B1(_1089_),
    .X(_1413_));
 sky130_fd_sc_hd__o21ai_1 _4331_ (.A1(_1226_),
    .A2(net30),
    .B1(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__nand2_1 _4332_ (.A(_1390_),
    .B(\datapath.RegB[7] ),
    .Y(_1415_));
 sky130_fd_sc_hd__a21oi_1 _4333_ (.A1(_1414_),
    .A2(_1415_),
    .B1(_1545_),
    .Y(_0050_));
 sky130_fd_sc_hd__a21o_1 _4334_ (.A1(\datapath.RegB[7] ),
    .A2(_1376_),
    .B1(_1089_),
    .X(_1416_));
 sky130_fd_sc_hd__o21ai_1 _4335_ (.A1(_1226_),
    .A2(net31),
    .B1(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__nand2_1 _4336_ (.A(_1390_),
    .B(\datapath.RegB[8] ),
    .Y(_1418_));
 sky130_fd_sc_hd__a21oi_1 _4337_ (.A1(_1417_),
    .A2(_1418_),
    .B1(_1545_),
    .Y(_0051_));
 sky130_fd_sc_hd__a21o_1 _4338_ (.A1(\datapath.RegB[8] ),
    .A2(_1376_),
    .B1(\control_unit.LoadA ),
    .X(_1420_));
 sky130_fd_sc_hd__o21ai_1 _4339_ (.A1(_1226_),
    .A2(net32),
    .B1(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__nand2_1 _4340_ (.A(_1390_),
    .B(\datapath.RegB[9] ),
    .Y(_1422_));
 sky130_fd_sc_hd__a21oi_1 _4341_ (.A1(_1421_),
    .A2(_1422_),
    .B1(_1545_),
    .Y(_0052_));
 sky130_fd_sc_hd__a21o_1 _4342_ (.A1(\datapath.RegB[9] ),
    .A2(_1376_),
    .B1(\control_unit.LoadA ),
    .X(_1423_));
 sky130_fd_sc_hd__o21ai_1 _4343_ (.A1(_1226_),
    .A2(net18),
    .B1(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__nand2_1 _4344_ (.A(_1390_),
    .B(\datapath.RegB[10] ),
    .Y(_1425_));
 sky130_fd_sc_hd__a21oi_1 _4345_ (.A1(_1424_),
    .A2(_1425_),
    .B1(_1544_),
    .Y(_0053_));
 sky130_fd_sc_hd__a21o_1 _4346_ (.A1(\datapath.RegB[10] ),
    .A2(_1376_),
    .B1(\control_unit.LoadA ),
    .X(_1426_));
 sky130_fd_sc_hd__o21ai_1 _4347_ (.A1(_1226_),
    .A2(net19),
    .B1(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__nand2_1 _4348_ (.A(_1390_),
    .B(\datapath.RegB[11] ),
    .Y(_1428_));
 sky130_fd_sc_hd__a21oi_1 _4349_ (.A1(_1427_),
    .A2(_1428_),
    .B1(_1544_),
    .Y(_0054_));
 sky130_fd_sc_hd__a21o_1 _4350_ (.A1(\datapath.RegB[11] ),
    .A2(_1376_),
    .B1(\control_unit.LoadA ),
    .X(_1429_));
 sky130_fd_sc_hd__o21ai_1 _4351_ (.A1(_1226_),
    .A2(net20),
    .B1(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__nand2_1 _4352_ (.A(_1390_),
    .B(\datapath.RegB[12] ),
    .Y(_1431_));
 sky130_fd_sc_hd__a21oi_1 _4353_ (.A1(_1430_),
    .A2(_1431_),
    .B1(_1544_),
    .Y(_0055_));
 sky130_fd_sc_hd__a21o_1 _4354_ (.A1(\datapath.RegB[12] ),
    .A2(_1376_),
    .B1(\control_unit.LoadA ),
    .X(_1432_));
 sky130_fd_sc_hd__o21ai_1 _4355_ (.A1(_1226_),
    .A2(net21),
    .B1(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__nand2_1 _4356_ (.A(_1390_),
    .B(\datapath.RegB[13] ),
    .Y(_1434_));
 sky130_fd_sc_hd__a21oi_1 _4357_ (.A1(_1433_),
    .A2(_1434_),
    .B1(_1544_),
    .Y(_0056_));
 sky130_fd_sc_hd__nand2_1 _4358_ (.A(_1390_),
    .B(\datapath.RegB[14] ),
    .Y(_1436_));
 sky130_fd_sc_hd__nand3_1 _4359_ (.A(_1045_),
    .B(\datapath.RegB[13] ),
    .C(_1376_),
    .Y(_1437_));
 sky130_fd_sc_hd__nand2_1 _4360_ (.A(_1089_),
    .B(net22),
    .Y(_1438_));
 sky130_fd_sc_hd__a31oi_1 _4361_ (.A1(_1436_),
    .A2(_1437_),
    .A3(_1438_),
    .B1(_1544_),
    .Y(_0057_));
 sky130_fd_sc_hd__and3_1 _4362_ (.A(_1045_),
    .B(\datapath.RegB[14] ),
    .C(_1376_),
    .X(_1439_));
 sky130_fd_sc_hd__a221o_1 _4363_ (.A1(_1089_),
    .A2(net23),
    .B1(\control_unit.regBk ),
    .B2(_1390_),
    .C1(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__nand2_1 _4364_ (.A(_1440_),
    .B(_1078_),
    .Y(_1441_));
 sky130_fd_sc_hd__clkinv_2 _4365_ (.A(_1441_),
    .Y(_0058_));
 sky130_fd_sc_hd__buf_1 _4366_ (.A(clknet_2_2__leaf_clk),
    .X(_1442_));
 sky130_fd_sc_hd__inv_2 _4368__2 (.A(clknet_1_0__leaf__1442_),
    .Y(net69));
 sky130_fd_sc_hd__inv_2 _4369__3 (.A(clknet_1_0__leaf__1442_),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _4370__4 (.A(clknet_1_0__leaf__1442_),
    .Y(net71));
 sky130_fd_sc_hd__inv_2 _4371__5 (.A(clknet_1_1__leaf__1442_),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _4372__6 (.A(clknet_1_1__leaf__1442_),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _4373__7 (.A(clknet_1_1__leaf__1442_),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _4374__8 (.A(clknet_1_1__leaf__1442_),
    .Y(net75));
 sky130_fd_sc_hd__inv_2 _4375__9 (.A(clknet_1_0__leaf__1442_),
    .Y(net76));
 sky130_fd_sc_hd__inv_2 _4376__10 (.A(clknet_1_0__leaf__1442_),
    .Y(net77));
 sky130_fd_sc_hd__inv_2 _4377__11 (.A(clknet_1_1__leaf__1442_),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _4378__12 (.A(clknet_1_1__leaf__1442_),
    .Y(net79));
 sky130_fd_sc_hd__inv_2 _4379__13 (.A(clknet_1_1__leaf__1442_),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _4380__14 (.A(clknet_1_0__leaf__1442_),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _4381__15 (.A(clknet_1_1__leaf__1442_),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _4382__16 (.A(clknet_1_1__leaf__1442_),
    .Y(net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__inv_2 _4383_ (.A(\control_unit.LoadCoun ),
    .Y(_1444_));
 sky130_fd_sc_hd__nor2_1 _4384_ (.A(\datapath.Counter[0] ),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__and2_1 _4385_ (.A(_1444_),
    .B(\datapath.Counter[0] ),
    .X(_1446_));
 sky130_fd_sc_hd__a211o_1 _4386_ (.A1(_1445_),
    .A2(\control_unit.S_Coun ),
    .B1(_1544_),
    .C1(_1446_),
    .X(_0075_));
 sky130_fd_sc_hd__or2_1 _4387_ (.A(\datapath.Counter[1] ),
    .B(_1445_),
    .X(_1447_));
 sky130_fd_sc_hd__o21a_1 _4388_ (.A1(\control_unit.S_Coun ),
    .A2(_1444_),
    .B1(_1067_),
    .X(_1449_));
 sky130_fd_sc_hd__nand2_1 _4389_ (.A(_1445_),
    .B(\datapath.Counter[1] ),
    .Y(_1450_));
 sky130_fd_sc_hd__and3_1 _4390_ (.A(_1447_),
    .B(_1449_),
    .C(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__clkbuf_1 _4391_ (.A(_1451_),
    .X(_0076_));
 sky130_fd_sc_hd__o31ai_1 _4392_ (.A1(\datapath.Counter[1] ),
    .A2(\datapath.Counter[0] ),
    .A3(_1444_),
    .B1(\datapath.Counter[2] ),
    .Y(_1452_));
 sky130_fd_sc_hd__nand2_1 _4393_ (.A(_1445_),
    .B(_1477_),
    .Y(_1453_));
 sky130_fd_sc_hd__inv_2 _4394_ (.A(_1449_),
    .Y(_1454_));
 sky130_fd_sc_hd__a21oi_1 _4395_ (.A1(_1452_),
    .A2(_1453_),
    .B1(_1454_),
    .Y(_0077_));
 sky130_fd_sc_hd__nor2_1 _4396_ (.A(\datapath.Counter[3] ),
    .B(_1453_),
    .Y(_1455_));
 sky130_fd_sc_hd__inv_2 _4397_ (.A(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__nand2_1 _4398_ (.A(_1453_),
    .B(\datapath.Counter[3] ),
    .Y(_1458_));
 sky130_fd_sc_hd__a21o_1 _4399_ (.A1(_1456_),
    .A2(_1458_),
    .B1(_1454_),
    .X(_1459_));
 sky130_fd_sc_hd__clkinv_2 _4400_ (.A(_1459_),
    .Y(_0078_));
 sky130_fd_sc_hd__or2_1 _4401_ (.A(\datapath.Counter[4] ),
    .B(_1455_),
    .X(_1460_));
 sky130_fd_sc_hd__nand2_1 _4402_ (.A(_1455_),
    .B(\datapath.Counter[4] ),
    .Y(_1461_));
 sky130_fd_sc_hd__a21o_1 _4403_ (.A1(_1460_),
    .A2(_1461_),
    .B1(_1454_),
    .X(_0079_));
 sky130_fd_sc_hd__dfxtp_1 _4404_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0016_),
    .Q(\datapath.MultiplierAC.PPG0.X[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4405_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0017_),
    .Q(\datapath.MultiplierAC.PPG0.X[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4406_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0018_),
    .Q(\datapath.MultiplierAC.PPG0.X[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4407_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0019_),
    .Q(\datapath.MultiplierAC.PPG0.X[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4408_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0020_),
    .Q(\datapath.MultiplierAC.PPG0.X[4] ));
 sky130_fd_sc_hd__dfxtp_4 _4409_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0021_),
    .Q(\datapath.MultiplierAC.PPG0.X[5] ));
 sky130_fd_sc_hd__dfxtp_2 _4410_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0022_),
    .Q(\datapath.MultiplierAC.PPG0.X[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4411_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0023_),
    .Q(\datapath.MultiplierAC.PPG0.X[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4412_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0024_),
    .Q(\datapath.MultiplierAC.PPG0.X[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4413_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0025_),
    .Q(\datapath.MultiplierAC.PPG0.X[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4414_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0026_),
    .Q(\datapath.MultiplierAC.PPG0.X[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4415_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0027_),
    .Q(\datapath.MultiplierAC.PPG0.X[11] ));
 sky130_fd_sc_hd__dfxtp_4 _4416_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0028_),
    .Q(\datapath.MultiplierAC.PPG0.X[12] ));
 sky130_fd_sc_hd__dfxtp_2 _4417_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0029_),
    .Q(\datapath.MultiplierAC.PPG0.X[13] ));
 sky130_fd_sc_hd__dfxtp_2 _4418_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0030_),
    .Q(\datapath.MultiplierAC.PPG0.X[14] ));
 sky130_fd_sc_hd__dfxtp_2 _4419_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0031_),
    .Q(\datapath.MultiplierAC.PPG0.X[15] ));
 sky130_fd_sc_hd__dfxtp_2 _4420_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0032_),
    .Q(\control_unit.S_C[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4421_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0033_),
    .Q(\control_unit.S_C[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4422_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0034_),
    .Q(\control_unit.S_Coun ));
 sky130_fd_sc_hd__dfxtp_1 _4423_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0035_),
    .Q(\control_unit.LoadC ));
 sky130_fd_sc_hd__dfxtp_1 _4424_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0036_),
    .Q(\control_unit.ShiftB ));
 sky130_fd_sc_hd__dfxtp_4 _4425_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0037_),
    .Q(\control_unit.LoadA ));
 sky130_fd_sc_hd__dfxtp_1 _4426_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0038_),
    .Q(\control_unit.LoadCoun ));
 sky130_fd_sc_hd__dfxtp_1 _4427_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0039_),
    .Q(\control_unit.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4428_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0040_),
    .Q(\control_unit.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4429_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0041_),
    .Q(\control_unit.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4430_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0042_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _4431_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0043_),
    .Q(\datapath.RegB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4432_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0044_),
    .Q(\datapath.RegB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4433_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0045_),
    .Q(\datapath.RegB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4434_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0046_),
    .Q(\datapath.RegB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4435_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0047_),
    .Q(\datapath.RegB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4436_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0048_),
    .Q(\datapath.RegB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4437_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0049_),
    .Q(\datapath.RegB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4438_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0050_),
    .Q(\datapath.RegB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4439_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0051_),
    .Q(\datapath.RegB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4440_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0052_),
    .Q(\datapath.RegB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4441_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0053_),
    .Q(\datapath.RegB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4442_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0054_),
    .Q(\datapath.RegB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4443_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0055_),
    .Q(\datapath.RegB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4444_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0056_),
    .Q(\datapath.RegB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4445_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0057_),
    .Q(\datapath.RegB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4446_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0058_),
    .Q(\control_unit.regBk ));
 sky130_fd_sc_hd__dfxtp_1 _4447_ (.CLK(net68),
    .D(_0059_),
    .Q(\datapath.MultiplierAC.PPG0.Y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4448_ (.CLK(net69),
    .D(_0060_),
    .Q(\datapath.MultiplierAC.PPG0.Y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4449_ (.CLK(net70),
    .D(_0061_),
    .Q(\datapath.MultiplierAC.PPG0.Y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4450_ (.CLK(net71),
    .D(_0062_),
    .Q(\datapath.MultiplierAC.PPG0.Y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4451_ (.CLK(net72),
    .D(_0063_),
    .Q(\datapath.MultiplierAC.PPG0.Y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4452_ (.CLK(net73),
    .D(_0064_),
    .Q(\datapath.MultiplierAC.PPG0.Y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4453_ (.CLK(net74),
    .D(_0065_),
    .Q(\datapath.MultiplierAC.PPG0.Y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4454_ (.CLK(net75),
    .D(_0066_),
    .Q(\datapath.MultiplierAC.PPG0.Y[7] ));
 sky130_fd_sc_hd__dfxtp_2 _4455_ (.CLK(net76),
    .D(_0067_),
    .Q(\datapath.MultiplierAC.PPG0.Y[8] ));
 sky130_fd_sc_hd__dfxtp_2 _4456_ (.CLK(net77),
    .D(_0068_),
    .Q(\datapath.MultiplierAC.PPG0.Y[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4457_ (.CLK(net78),
    .D(_0069_),
    .Q(\datapath.MultiplierAC.PPG0.Y[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4458_ (.CLK(net79),
    .D(_0070_),
    .Q(\datapath.MultiplierAC.PPG0.Y[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4459_ (.CLK(net80),
    .D(_0071_),
    .Q(\datapath.MultiplierAC.PPG0.Y[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4460_ (.CLK(net81),
    .D(_0072_),
    .Q(\datapath.MultiplierAC.PPG0.Y[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4461_ (.CLK(net82),
    .D(_0073_),
    .Q(\datapath.MultiplierAC.PPG0.Y[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4462_ (.CLK(net83),
    .D(_0074_),
    .Q(\datapath.MultiplierAC.PPG0.Y[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4463_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0075_),
    .Q(\datapath.Counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4464_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0076_),
    .Q(\datapath.Counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4465_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0077_),
    .Q(\datapath.Counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4466_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0078_),
    .Q(\datapath.Counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4467_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0079_),
    .Q(\datapath.Counter[4] ));
 sky130_fd_sc_hd__conb_1 L2RExp_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 L2RExp_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 L2RExp_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 L2RExp_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 L2RExp_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 L2RExp_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 L2RExp_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 L2RExp_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 L2RExp_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 L2RExp_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 L2RExp_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 L2RExp_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 L2RExp_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 L2RExp_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 L2RExp_67 (.LO(net67));
 sky130_fd_sc_hd__inv_2 _4367__1 (.A(clknet_1_0__leaf__1442_),
    .Y(net68));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(A[1]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(A[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(A[3]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(A[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(A[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(A[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(A[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(A[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(A[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(B[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(B[10]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(B[11]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(B[12]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(B[13]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(B[14]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(B[15]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(B[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(B[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(B[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(B[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(B[5]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(B[6]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(B[7]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(B[8]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(B[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(rst),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(start),
    .X(net34));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(C[0]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(C[10]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(C[11]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(C[12]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(C[13]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(C[14]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(C[15]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(C[1]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(C[2]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(C[3]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(C[4]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(C[5]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(C[6]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(C[7]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(C[8]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(C[9]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(Done));
 sky130_fd_sc_hd__conb_1 L2RExp_52 (.LO(net52));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1442_ (.A(_1442_),
    .X(clknet_0__1442_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1442_ (.A(clknet_0__1442_),
    .X(clknet_1_0__leaf__1442_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1442_ (.A(clknet_0__1442_),
    .X(clknet_1_1__leaf__1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net24));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_405 ();
 assign C[16] = net52;
 assign C[17] = net53;
 assign C[18] = net54;
 assign C[19] = net55;
 assign C[20] = net56;
 assign C[21] = net57;
 assign C[22] = net58;
 assign C[23] = net59;
 assign C[24] = net60;
 assign C[25] = net61;
 assign C[26] = net62;
 assign C[27] = net63;
 assign C[28] = net64;
 assign C[29] = net65;
 assign C[30] = net66;
 assign C[31] = net67;
endmodule
